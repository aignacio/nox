`ifndef _NOX_UTILS_PKG_
`define _NOX_UTILS_PKG_
  package nox_utils_pkg;
    `include "nox_pkg.svh"
    `include "core_bus_pkg.svh"
    `include "riscv_pkg.svh"
  endpackage
`endif
