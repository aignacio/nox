module boot_rom (
  input          clk,
  input          en,
  input  [12:0]  addr_i,
  output [31:0]  dout_o
);

 // Based on this UG - https://www.xilinx.com/support/documentation/sw_manuals/xilinx2020_1/ug901-vivado-synthesis.pdf

 (*rom_style = "block" *) logic [31:0] data;
 assign dout_o = data;

 always @(posedge clk) begin
     if (en) begin
         case (addr_i)
         'd0: data <= 32'h90001197;         'd1: data <= 32'h80018193;
         'd2: data <= 32'h90002117;         'd3: data <= 32'hff810113;
         'd4: data <= 32'h004000ef;         'd5: data <= 32'h800007b7;
         'd6: data <= 32'h10178793;         'd7: data <= 32'h30579073;
         'd8: data <= 32'h800067b7;         'd9: data <= 32'h84478493;
         'd10: data <= 32'h100007b7;         'd11: data <= 32'h00078093;
         'd12: data <= 32'h0140006f;         'd13: data <= 32'h0004a783;
         'd14: data <= 32'h00f0a023;         'd15: data <= 32'h00408093;
         'd16: data <= 32'h00448493;         'd17: data <= 32'h87818793;
         'd18: data <= 32'hfef0e6e3;         'd19: data <= 32'h87818093;
         'd20: data <= 32'h00c0006f;         'd21: data <= 32'h0000a023;
         'd22: data <= 32'h00408093;         'd23: data <= 32'h89018793;
         'd24: data <= 32'hfef0eae3;         'd25: data <= 32'h7f5000ef;
         'd26: data <= 32'h00000013;         'd27: data <= 32'h00000000;
         'd28: data <= 32'h00000000;         'd29: data <= 32'h00000000;
         'd30: data <= 32'h00000000;         'd31: data <= 32'h00000000;
         'd32: data <= 32'h00000000;         'd33: data <= 32'h00000000;
         'd34: data <= 32'h00000000;         'd35: data <= 32'h00000000;
         'd36: data <= 32'h00000000;         'd37: data <= 32'h00000000;
         'd38: data <= 32'h00000000;         'd39: data <= 32'h00000000;
         'd40: data <= 32'h00000000;         'd41: data <= 32'h00000000;
         'd42: data <= 32'h00000000;         'd43: data <= 32'h00000000;
         'd44: data <= 32'h00000000;         'd45: data <= 32'h00000000;
         'd46: data <= 32'h00000000;         'd47: data <= 32'h00000000;
         'd48: data <= 32'h00000000;         'd49: data <= 32'h00000000;
         'd50: data <= 32'h00000000;         'd51: data <= 32'h00000000;
         'd52: data <= 32'h00000000;         'd53: data <= 32'h00000000;
         'd54: data <= 32'h00000000;         'd55: data <= 32'h00000000;
         'd56: data <= 32'h00000000;         'd57: data <= 32'h00000000;
         'd58: data <= 32'h00000000;         'd59: data <= 32'h00000000;
         'd60: data <= 32'h00000000;         'd61: data <= 32'h00000000;
         'd62: data <= 32'h00000000;         'd63: data <= 32'h00000000;
         'd64: data <= 32'hfd010113;         'd65: data <= 32'h02112623;
         'd66: data <= 32'h02812423;         'd67: data <= 32'h03010413;
         'd68: data <= 32'hfca42e23;         'd69: data <= 32'hfcb42c23;
         'd70: data <= 32'hfdc42783;         'd71: data <= 32'h0007d783;
         'd72: data <= 32'hfef41523;         'd73: data <= 32'hfea41783;
         'd74: data <= 32'h4077d793;         'd75: data <= 32'h01079793;
         'd76: data <= 32'h4107d793;         'd77: data <= 32'h0ff7f793;
         'd78: data <= 32'h0017f793;         'd79: data <= 32'hfef404a3;
         'd80: data <= 32'hfe944783;         'd81: data <= 32'h00078c63;
         'd82: data <= 32'hfea45783;         'd83: data <= 32'h07f7f793;
         'd84: data <= 32'h01079793;         'd85: data <= 32'h4107d793;
         'd86: data <= 32'h18c0006f;         'd87: data <= 32'hfea45783;
         'd88: data <= 32'h0077f793;         'd89: data <= 32'hfef41323;
         'd90: data <= 32'hfea41783;         'd91: data <= 32'h4037d793;
         'd92: data <= 32'h01079793;         'd93: data <= 32'h4107d793;
         'd94: data <= 32'h00f7f793;         'd95: data <= 32'hfef41623;
         'd96: data <= 32'hfec41783;         'd97: data <= 32'h00479793;
         'd98: data <= 32'h01079713;         'd99: data <= 32'h41075713;
         'd100: data <= 32'hfec45783;         'd101: data <= 32'h00f767b3;
         'd102: data <= 32'hfef41623;         'd103: data <= 32'hfe641783;
         'd104: data <= 32'h00078863;         'd105: data <= 32'h00100713;
         'd106: data <= 32'h06e78863;         'd107: data <= 32'h0b40006f;
         'd108: data <= 32'hfec41703;         'd109: data <= 32'h02100793;
         'd110: data <= 32'h00e7c663;         'd111: data <= 32'h02200793;
         'd112: data <= 32'hfef41623;         'd113: data <= 32'hfd842783;
         'd114: data <= 32'h0187a503;         'd115: data <= 32'hfd842783;
         'd116: data <= 32'h0147a583;         'd117: data <= 32'hfd842783;
         'd118: data <= 32'h00079603;         'd119: data <= 32'hfd842783;
         'd120: data <= 32'h00279683;         'd121: data <= 32'hfd842783;
         'd122: data <= 32'h0387d783;         'd123: data <= 32'hfec41703;
         'd124: data <= 32'h1dd020ef;         'd125: data <= 32'h00050793;
         'd126: data <= 32'hfef41723;         'd127: data <= 32'hfd842783;
         'd128: data <= 32'h03e7d783;         'd129: data <= 32'h06079463;
         'd130: data <= 32'hfee45703;         'd131: data <= 32'hfd842783;
         'd132: data <= 32'h02e79f23;         'd133: data <= 32'h0580006f;
         'd134: data <= 32'hfd842783;         'd135: data <= 32'h02878713;
         'd136: data <= 32'hfd842783;         'd137: data <= 32'h0387d683;
         'd138: data <= 32'hfec41783;         'd139: data <= 32'h00068613;
         'd140: data <= 32'h00078593;         'd141: data <= 32'h00070513;
         'd142: data <= 32'h531010ef;         'd143: data <= 32'h00050793;
         'd144: data <= 32'hfef41723;         'd145: data <= 32'hfd842783;
         'd146: data <= 32'h03c7d783;         'd147: data <= 32'h02079463;
         'd148: data <= 32'hfee45703;         'd149: data <= 32'hfd842783;
         'd150: data <= 32'h02e79e23;         'd151: data <= 32'h0180006f;
         'd152: data <= 32'hfea45783;         'd153: data <= 32'hfef41723;
         'd154: data <= 32'h0100006f;         'd155: data <= 32'h00000013;
         'd156: data <= 32'h0080006f;         'd157: data <= 32'h00000013;
         'd158: data <= 32'hfee45703;         'd159: data <= 32'hfd842783;
         'd160: data <= 32'h0387d783;         'd161: data <= 32'h00078593;
         'd162: data <= 32'h00070513;         'd163: data <= 32'h3e0030ef;
         'd164: data <= 32'h00050793;         'd165: data <= 32'h00078713;
         'd166: data <= 32'hfd842783;         'd167: data <= 32'h02e79c23;
         'd168: data <= 32'hfee45783;         'd169: data <= 32'h07f7f793;
         'd170: data <= 32'hfef41723;         'd171: data <= 32'hfea45783;
         'd172: data <= 32'hf007f793;         'd173: data <= 32'h01079793;
         'd174: data <= 32'h4107d793;         'd175: data <= 32'h0807e793;
         'd176: data <= 32'h01079713;         'd177: data <= 32'h41075713;
         'd178: data <= 32'hfee45783;         'd179: data <= 32'h00f767b3;
         'd180: data <= 32'h01079713;         'd181: data <= 32'h41075713;
         'd182: data <= 32'hfdc42783;         'd183: data <= 32'h00e79023;
         'd184: data <= 32'hfee41783;         'd185: data <= 32'h00078513;
         'd186: data <= 32'h02c12083;         'd187: data <= 32'h02812403;
         'd188: data <= 32'h03010113;         'd189: data <= 32'h00008067;
         'd190: data <= 32'hfd010113;         'd191: data <= 32'h02112623;
         'd192: data <= 32'h02812423;         'd193: data <= 32'h03010413;
         'd194: data <= 32'hfca42e23;         'd195: data <= 32'hfcb42c23;
         'd196: data <= 32'hfcc42a23;         'd197: data <= 32'hfdc42783;
         'd198: data <= 32'hfd442583;         'd199: data <= 32'h00078513;
         'd200: data <= 32'hde1ff0ef;         'd201: data <= 32'h00050793;
         'd202: data <= 32'hfef41723;         'd203: data <= 32'hfd842783;
         'd204: data <= 32'hfd442583;         'd205: data <= 32'h00078513;
         'd206: data <= 32'hdc9ff0ef;         'd207: data <= 32'h00050793;
         'd208: data <= 32'hfef41623;         'd209: data <= 32'hfee41703;
         'd210: data <= 32'hfec41783;         'd211: data <= 32'h40f707b3;
         'd212: data <= 32'h00078513;         'd213: data <= 32'h02c12083;
         'd214: data <= 32'h02812403;         'd215: data <= 32'h03010113;
         'd216: data <= 32'h00008067;         'd217: data <= 32'hfe010113;
         'd218: data <= 32'h00812e23;         'd219: data <= 32'h02010413;
         'd220: data <= 32'hfea42623;         'd221: data <= 32'hfeb42423;
         'd222: data <= 32'hfec42223;         'd223: data <= 32'hfe442783;
         'd224: data <= 32'h08079e63;         'd225: data <= 32'hfec42783;
         'd226: data <= 32'h00079783;         'd227: data <= 32'hf007f793;
         'd228: data <= 32'h01079713;         'd229: data <= 32'h41075713;
         'd230: data <= 32'hfec42783;         'd231: data <= 32'h00079783;
         'd232: data <= 32'h01079793;         'd233: data <= 32'h0107d793;
         'd234: data <= 32'h0087d793;         'd235: data <= 32'h01079793;
         'd236: data <= 32'h0107d793;         'd237: data <= 32'h01079793;
         'd238: data <= 32'h4107d793;         'd239: data <= 32'h00f767b3;
         'd240: data <= 32'h01079713;         'd241: data <= 32'h41075713;
         'd242: data <= 32'hfec42783;         'd243: data <= 32'h00e79023;
         'd244: data <= 32'hfe842783;         'd245: data <= 32'h00079783;
         'd246: data <= 32'hf007f793;         'd247: data <= 32'h01079713;
         'd248: data <= 32'h41075713;         'd249: data <= 32'hfe842783;
         'd250: data <= 32'h00079783;         'd251: data <= 32'h01079793;
         'd252: data <= 32'h0107d793;         'd253: data <= 32'h0087d793;
         'd254: data <= 32'h01079793;         'd255: data <= 32'h0107d793;
         'd256: data <= 32'h01079793;         'd257: data <= 32'h4107d793;
         'd258: data <= 32'h00f767b3;         'd259: data <= 32'h01079713;
         'd260: data <= 32'h41075713;         'd261: data <= 32'hfe842783;
         'd262: data <= 32'h00e79023;         'd263: data <= 32'hfec42783;
         'd264: data <= 32'h00279783;         'd265: data <= 32'h00078713;
         'd266: data <= 32'hfe842783;         'd267: data <= 32'h00279783;
         'd268: data <= 32'h40f707b3;         'd269: data <= 32'h00078513;
         'd270: data <= 32'h01c12403;         'd271: data <= 32'h02010113;
         'd272: data <= 32'h00008067;         'd273: data <= 32'hfe010113;
         'd274: data <= 32'h00812e23;         'd275: data <= 32'h02010413;
         'd276: data <= 32'hfea42623;         'd277: data <= 32'hfeb42423;
         'd278: data <= 32'hfe842783;         'd279: data <= 32'h00079703;
         'd280: data <= 32'hfec42783;         'd281: data <= 32'h00e79023;
         'd282: data <= 32'hfe842783;         'd283: data <= 32'h00279703;
         'd284: data <= 32'hfec42783;         'd285: data <= 32'h00e79123;
         'd286: data <= 32'h00000013;         'd287: data <= 32'h01c12403;
         'd288: data <= 32'h02010113;         'd289: data <= 32'h00008067;
         'd290: data <= 32'hfc010113;         'd291: data <= 32'h02112e23;
         'd292: data <= 32'h02812c23;         'd293: data <= 32'h04010413;
         'd294: data <= 32'hfca42623;         'd295: data <= 32'h00058793;
         'd296: data <= 32'hfcf41523;         'd297: data <= 32'hfe041723;
         'd298: data <= 32'hfe041623;         'd299: data <= 32'hfe041523;
         'd300: data <= 32'hfcc42783;         'd301: data <= 32'h0247a783;
         'd302: data <= 32'hfef42223;         'd303: data <= 32'hfcc42783;
         'd304: data <= 32'h0047d783;         'd305: data <= 32'hfcf41e23;
         'd306: data <= 32'hfca45783;         'd307: data <= 32'hfcf41923;
         'd308: data <= 32'hfc041f23;         'd309: data <= 32'h1780006f;
         'd310: data <= 32'hfde45783;         'd311: data <= 32'h0ff7f793;
         'd312: data <= 32'h01079793;         'd313: data <= 32'h4107d793;
         'd314: data <= 32'hfcf41823;         'd315: data <= 32'hfd040793;
         'd316: data <= 32'h00078593;         'd317: data <= 32'hfe442503;
         'd318: data <= 32'h748000ef;         'd319: data <= 32'hfca42a23;
         'd320: data <= 32'hfe442503;         'd321: data <= 32'h7e0000ef;
         'd322: data <= 32'hfea42223;         'd323: data <= 32'hfd442783;
         'd324: data <= 32'h04079863;         'd325: data <= 32'hfea45783;
         'd326: data <= 32'h00178793;         'd327: data <= 32'hfef41523;
         'd328: data <= 32'hfe442783;         'd329: data <= 32'h0007a783;
         'd330: data <= 32'h0047a783;         'd331: data <= 32'h00079783;
         'd332: data <= 32'h4087d793;         'd333: data <= 32'h01079793;
         'd334: data <= 32'h4107d793;         'd335: data <= 32'h01079793;
         'd336: data <= 32'h0107d793;         'd337: data <= 32'h0017f793;
         'd338: data <= 32'h01079713;         'd339: data <= 32'h01075713;
         'd340: data <= 32'hfee45783;         'd341: data <= 32'h00f707b3;
         'd342: data <= 32'hfef41723;         'd343: data <= 32'h0a80006f;
         'd344: data <= 32'hfec45783;         'd345: data <= 32'h00178793;
         'd346: data <= 32'hfef41623;         'd347: data <= 32'hfd442783;
         'd348: data <= 32'h0047a783;         'd349: data <= 32'h00079783;
         'd350: data <= 32'h01079793;         'd351: data <= 32'h0107d793;
         'd352: data <= 32'h0017f793;         'd353: data <= 32'h02078e63;
         'd354: data <= 32'hfd442783;         'd355: data <= 32'h0047a783;
         'd356: data <= 32'h00079783;         'd357: data <= 32'h4097d793;
         'd358: data <= 32'h01079793;         'd359: data <= 32'h4107d793;
         'd360: data <= 32'h01079793;         'd361: data <= 32'h0107d793;
         'd362: data <= 32'h0017f793;         'd363: data <= 32'h01079713;
         'd364: data <= 32'h01075713;         'd365: data <= 32'hfee45783;
         'd366: data <= 32'h00f707b3;         'd367: data <= 32'hfef41723;
         'd368: data <= 32'hfd442783;         'd369: data <= 32'h0007a783;
         'd370: data <= 32'h02078e63;         'd371: data <= 32'hfd442783;
         'd372: data <= 32'h0007a783;         'd373: data <= 32'hfef42023;
         'd374: data <= 32'hfe042783;         'd375: data <= 32'h0007a703;
         'd376: data <= 32'hfd442783;         'd377: data <= 32'h00e7a023;
         'd378: data <= 32'hfe442783;         'd379: data <= 32'h0007a703;
         'd380: data <= 32'hfe042783;         'd381: data <= 32'h00e7a023;
         'd382: data <= 32'hfe442783;         'd383: data <= 32'hfe042703;
         'd384: data <= 32'h00e7a023;         'd385: data <= 32'hfd241783;
         'd386: data <= 32'h0207c463;         'd387: data <= 32'hfd241783;
         'd388: data <= 32'h01079793;         'd389: data <= 32'h0107d793;
         'd390: data <= 32'h00178793;         'd391: data <= 32'h01079793;
         'd392: data <= 32'h0107d793;         'd393: data <= 32'h01079793;
         'd394: data <= 32'h4107d793;         'd395: data <= 32'hfcf41923;
         'd396: data <= 32'hfde41783;         'd397: data <= 32'h01079793;
         'd398: data <= 32'h0107d793;         'd399: data <= 32'h00178793;
         'd400: data <= 32'h01079793;         'd401: data <= 32'h0107d793;
         'd402: data <= 32'hfcf41f23;         'd403: data <= 32'hfde41703;
         'd404: data <= 32'hfdc41783;         'd405: data <= 32'he8f742e3;
         'd406: data <= 32'hfec45783;         'd407: data <= 32'h00279793;
         'd408: data <= 32'h01079713;         'd409: data <= 32'h01075713;
         'd410: data <= 32'hfea45783;         'd411: data <= 32'h40f707b3;
         'd412: data <= 32'h01079713;         'd413: data <= 32'h01075713;
         'd414: data <= 32'hfee45783;         'd415: data <= 32'h00f707b3;
         'd416: data <= 32'hfef41723;         'd417: data <= 32'hfca41783;
         'd418: data <= 32'h00f05e63;         'd419: data <= 32'hfcc42603;
         'd420: data <= 32'h800007b7;         'd421: data <= 32'h2f878593;
         'd422: data <= 32'hfe442503;         'd423: data <= 32'h6a4000ef;
         'd424: data <= 32'hfea42223;         'd425: data <= 32'hfe442783;
         'd426: data <= 32'h0007a783;         'd427: data <= 32'h00078513;
         'd428: data <= 32'h4b0000ef;         'd429: data <= 32'hfca42c23;
         'd430: data <= 32'hfd040793;         'd431: data <= 32'h00078593;
         'd432: data <= 32'hfe442503;         'd433: data <= 32'h57c000ef;
         'd434: data <= 32'hfea42023;         'd435: data <= 32'hfe042783;
         'd436: data <= 32'h04079263;         'd437: data <= 32'hfe442783;
         'd438: data <= 32'h0007a783;         'd439: data <= 32'hfef42023;
         'd440: data <= 32'h0340006f;         'd441: data <= 32'hfe442783;
         'd442: data <= 32'h0047a783;         'd443: data <= 32'h00079783;
         'd444: data <= 32'hfee45703;         'd445: data <= 32'h00070593;
         'd446: data <= 32'h00078513;         'd447: data <= 32'h078030ef;
         'd448: data <= 32'h00050793;         'd449: data <= 32'hfef41723;
         'd450: data <= 32'hfe042783;         'd451: data <= 32'h0007a783;
         'd452: data <= 32'hfef42023;         'd453: data <= 32'hfe042783;
         'd454: data <= 32'hfc0796e3;         'd455: data <= 32'hfe442783;
         'd456: data <= 32'h0007a783;         'd457: data <= 32'h00078593;
         'd458: data <= 32'hfd842503;         'd459: data <= 32'h4a8000ef;
         'd460: data <= 32'hfca42c23;         'd461: data <= 32'h00000613;
         'd462: data <= 32'h800007b7;         'd463: data <= 32'h36478593;
         'd464: data <= 32'hfe442503;         'd465: data <= 32'h5fc000ef;
         'd466: data <= 32'hfea42223;         'd467: data <= 32'hfe442783;
         'd468: data <= 32'h0007a783;         'd469: data <= 32'hfef42023;
         'd470: data <= 32'h0340006f;         'd471: data <= 32'hfe442783;
         'd472: data <= 32'h0047a783;         'd473: data <= 32'h00079783;
         'd474: data <= 32'hfee45703;         'd475: data <= 32'h00070593;
         'd476: data <= 32'h00078513;         'd477: data <= 32'h000030ef;
         'd478: data <= 32'h00050793;         'd479: data <= 32'hfef41723;
         'd480: data <= 32'hfe042783;         'd481: data <= 32'h0007a783;
         'd482: data <= 32'hfef42023;         'd483: data <= 32'hfe042783;
         'd484: data <= 32'hfc0796e3;         'd485: data <= 32'hfee45783;
         'd486: data <= 32'h00078513;         'd487: data <= 32'h03c12083;
         'd488: data <= 32'h03812403;         'd489: data <= 32'h04010113;
         'd490: data <= 32'h00008067;         'd491: data <= 32'hfb010113;
         'd492: data <= 32'h04112623;         'd493: data <= 32'h04812423;
         'd494: data <= 32'h05010413;         'd495: data <= 32'hfaa42e23;
         'd496: data <= 32'hfab42c23;         'd497: data <= 32'h00060793;
         'd498: data <= 32'hfaf41b23;         'd499: data <= 32'h01400793;
         'd500: data <= 32'hfef42223;         'd501: data <= 32'hfe442583;
         'd502: data <= 32'hfbc42503;         'd503: data <= 32'h77c040ef;
         'd504: data <= 32'h00050793;         'd505: data <= 32'hffe78793;
         'd506: data <= 32'hfef42023;         'd507: data <= 32'hfb842703;
         'd508: data <= 32'hfe042783;         'd509: data <= 32'h00379793;
         'd510: data <= 32'h00f707b3;         'd511: data <= 32'hfcf42e23;
         'd512: data <= 32'hfdc42783;         'd513: data <= 32'hfcf42423;
         'd514: data <= 32'hfc842703;         'd515: data <= 32'hfe042783;
         'd516: data <= 32'h00279793;         'd517: data <= 32'h00f707b3;
         'd518: data <= 32'hfcf42c23;         'd519: data <= 32'hfb842783;
         'd520: data <= 32'hfcf42a23;         'd521: data <= 32'hfd442783;
         'd522: data <= 32'h0007a023;         'd523: data <= 32'hfc842703;
         'd524: data <= 32'hfd442783;         'd525: data <= 32'h00e7a223;
         'd526: data <= 32'hfd442783;         'd527: data <= 32'h0047a783;
         'd528: data <= 32'h00079123;         'd529: data <= 32'hfd442783;
         'd530: data <= 32'h0047a783;         'd531: data <= 32'hffff8737;
         'd532: data <= 32'h08070713;         'd533: data <= 32'h00e79023;
         'd534: data <= 32'hfb842783;         'd535: data <= 32'h00878793;
         'd536: data <= 32'hfaf42c23;         'd537: data <= 32'hfc842783;
         'd538: data <= 32'h00478793;         'd539: data <= 32'hfcf42423;
         'd540: data <= 32'hffff87b7;         'd541: data <= 32'hfff7c793;
         'd542: data <= 32'hfcf41323;         'd543: data <= 32'hfff00793;
         'd544: data <= 32'hfcf41223;         'd545: data <= 32'hfc840693;
         'd546: data <= 32'hfb840613;         'd547: data <= 32'hfc440593;
         'd548: data <= 32'hfd842783;         'd549: data <= 32'hfdc42703;
         'd550: data <= 32'hfd442503;         'd551: data <= 32'h1d8000ef;
         'd552: data <= 32'hfe042623;         'd553: data <= 32'h0a40006f;
         'd554: data <= 32'hfec42783;         'd555: data <= 32'h01079713;
         'd556: data <= 32'h01075713;         'd557: data <= 32'hfb645783;
         'd558: data <= 32'h00f747b3;         'd559: data <= 32'h01079793;
         'd560: data <= 32'h0107d793;         'd561: data <= 32'h00f7f793;
         'd562: data <= 32'hfcf41823;         'd563: data <= 32'hfd045783;
         'd564: data <= 32'h00379793;         'd565: data <= 32'h01079713;
         'd566: data <= 32'h01075713;         'd567: data <= 32'hfec42783;
         'd568: data <= 32'h01079793;         'd569: data <= 32'h0107d793;
         'd570: data <= 32'h0077f793;         'd571: data <= 32'h01079793;
         'd572: data <= 32'h0107d793;         'd573: data <= 32'h00f767b3;
         'd574: data <= 32'hfcf41723;         'd575: data <= 32'hfce45783;
         'd576: data <= 32'h00879793;         'd577: data <= 32'h01079713;
         'd578: data <= 32'h41075713;         'd579: data <= 32'hfce41783;
         'd580: data <= 32'h00f767b3;         'd581: data <= 32'h01079793;
         'd582: data <= 32'h4107d793;         'd583: data <= 32'hfcf41223;
         'd584: data <= 32'hfc840693;         'd585: data <= 32'hfb840613;
         'd586: data <= 32'hfc440593;         'd587: data <= 32'hfd842783;
         'd588: data <= 32'hfdc42703;         'd589: data <= 32'hfd442503;
         'd590: data <= 32'h13c000ef;         'd591: data <= 32'hfec42783;
         'd592: data <= 32'h00178793;         'd593: data <= 32'hfef42623;
         'd594: data <= 32'hfec42703;         'd595: data <= 32'hfe042783;
         'd596: data <= 32'hf4f76ce3;         'd597: data <= 32'hfd442783;
         'd598: data <= 32'h0007a783;         'd599: data <= 32'hfef42423;
         'd600: data <= 32'h00100793;         'd601: data <= 32'hfef42623;
         'd602: data <= 32'h0d00006f;         'd603: data <= 32'hfe042783;
         'd604: data <= 32'h00500593;         'd605: data <= 32'h00078513;
         'd606: data <= 32'h5e0040ef;         'd607: data <= 32'h00050793;
         'd608: data <= 32'h00078713;         'd609: data <= 32'hfec42783;
         'd610: data <= 32'h02e7f463;         'd611: data <= 32'hfec42783;
         'd612: data <= 32'h00178713;         'd613: data <= 32'hfee42623;
         'd614: data <= 32'hfe842703;         'd615: data <= 32'h00472703;
         'd616: data <= 32'h01079793;         'd617: data <= 32'h4107d793;
         'd618: data <= 32'h00f71123;         'd619: data <= 32'h0800006f;
         'd620: data <= 32'hfec42783;         'd621: data <= 32'h00178713;
         'd622: data <= 32'hfee42623;         'd623: data <= 32'h01079713;
         'd624: data <= 32'h01075713;         'd625: data <= 32'hfb645783;
         'd626: data <= 32'h00f747b3;         'd627: data <= 32'hfcf41923;
         'd628: data <= 32'hfec42783;         'd629: data <= 32'h01079793;
         'd630: data <= 32'h0107d793;         'd631: data <= 32'h00879793;
         'd632: data <= 32'h01079793;         'd633: data <= 32'h0107d793;
         'd634: data <= 32'h7007f793;         'd635: data <= 32'h01079713;
         'd636: data <= 32'h01075713;         'd637: data <= 32'hfd245783;
         'd638: data <= 32'h00f767b3;         'd639: data <= 32'h01079793;
         'd640: data <= 32'h0107d793;         'd641: data <= 32'h01079693;
         'd642: data <= 32'h4106d693;         'd643: data <= 32'hfe842783;
         'd644: data <= 32'h0047a783;         'd645: data <= 32'h00004737;
         'd646: data <= 32'hfff70713;         'd647: data <= 32'h00e6f733;
         'd648: data <= 32'h01071713;         'd649: data <= 32'h41075713;
         'd650: data <= 32'h00e79123;         'd651: data <= 32'hfe842783;
         'd652: data <= 32'h0007a783;         'd653: data <= 32'hfef42423;
         'd654: data <= 32'hfe842783;         'd655: data <= 32'h0007a783;
         'd656: data <= 32'hf20796e3;         'd657: data <= 32'h00000613;
         'd658: data <= 32'h800007b7;         'd659: data <= 32'h36478593;
         'd660: data <= 32'hfd442503;         'd661: data <= 32'h2ec000ef;
         'd662: data <= 32'hfca42a23;         'd663: data <= 32'hfd442783;
         'd664: data <= 32'h00078513;         'd665: data <= 32'h04c12083;
         'd666: data <= 32'h04812403;         'd667: data <= 32'h05010113;
         'd668: data <= 32'h00008067;         'd669: data <= 32'hfc010113;
         'd670: data <= 32'h02112e23;         'd671: data <= 32'h02812c23;
         'd672: data <= 32'h04010413;         'd673: data <= 32'hfca42e23;
         'd674: data <= 32'hfcb42c23;         'd675: data <= 32'hfcc42a23;
         'd676: data <= 32'hfcd42823;         'd677: data <= 32'hfce42623;
         'd678: data <= 32'hfcf42423;         'd679: data <= 32'hfd442783;
         'd680: data <= 32'h0007a783;         'd681: data <= 32'h00878793;
         'd682: data <= 32'hfcc42703;         'd683: data <= 32'h00e7e663;
         'd684: data <= 32'h00000793;         'd685: data <= 32'h0980006f;
         'd686: data <= 32'hfd042783;         'd687: data <= 32'h0007a783;
         'd688: data <= 32'h00478793;         'd689: data <= 32'hfc842703;
         'd690: data <= 32'h00e7e663;         'd691: data <= 32'h00000793;
         'd692: data <= 32'h07c0006f;         'd693: data <= 32'hfd442783;
         'd694: data <= 32'h0007a783;         'd695: data <= 32'hfef42623;
         'd696: data <= 32'hfd442783;         'd697: data <= 32'h0007a783;
         'd698: data <= 32'h00878713;         'd699: data <= 32'hfd442783;
         'd700: data <= 32'h00e7a023;         'd701: data <= 32'hfdc42783;
         'd702: data <= 32'h0007a703;         'd703: data <= 32'hfec42783;
         'd704: data <= 32'h00e7a023;         'd705: data <= 32'hfdc42783;
         'd706: data <= 32'hfec42703;         'd707: data <= 32'h00e7a023;
         'd708: data <= 32'hfd042783;         'd709: data <= 32'h0007a703;
         'd710: data <= 32'hfec42783;         'd711: data <= 32'h00e7a223;
         'd712: data <= 32'hfd042783;         'd713: data <= 32'h0007a783;
         'd714: data <= 32'h00478713;         'd715: data <= 32'hfd042783;
         'd716: data <= 32'h00e7a023;         'd717: data <= 32'hfec42783;
         'd718: data <= 32'h0047a783;         'd719: data <= 32'hfd842583;
         'd720: data <= 32'h00078513;         'd721: data <= 32'h901ff0ef;
         'd722: data <= 32'hfec42783;         'd723: data <= 32'h00078513;
         'd724: data <= 32'h03c12083;         'd725: data <= 32'h03812403;
         'd726: data <= 32'h04010113;         'd727: data <= 32'h00008067;
         'd728: data <= 32'hfd010113;         'd729: data <= 32'h02812623;
         'd730: data <= 32'h03010413;         'd731: data <= 32'hfca42e23;
         'd732: data <= 32'hfdc42783;         'd733: data <= 32'h0007a783;
         'd734: data <= 32'hfef42623;         'd735: data <= 32'hfdc42783;
         'd736: data <= 32'h0047a783;         'd737: data <= 32'hfef42423;
         'd738: data <= 32'hfec42783;         'd739: data <= 32'h0047a703;
         'd740: data <= 32'hfdc42783;         'd741: data <= 32'h00e7a223;
         'd742: data <= 32'hfec42783;         'd743: data <= 32'hfe842703;
         'd744: data <= 32'h00e7a223;         'd745: data <= 32'hfdc42783;
         'd746: data <= 32'h0007a783;         'd747: data <= 32'h0007a703;
         'd748: data <= 32'hfdc42783;         'd749: data <= 32'h00e7a023;
         'd750: data <= 32'hfec42783;         'd751: data <= 32'h0007a023;
         'd752: data <= 32'hfec42783;         'd753: data <= 32'h00078513;
         'd754: data <= 32'h02c12403;         'd755: data <= 32'h03010113;
         'd756: data <= 32'h00008067;         'd757: data <= 32'hfd010113;
         'd758: data <= 32'h02812623;         'd759: data <= 32'h03010413;
         'd760: data <= 32'hfca42e23;         'd761: data <= 32'hfcb42c23;
         'd762: data <= 32'hfdc42783;         'd763: data <= 32'h0047a783;
         'd764: data <= 32'hfef42623;         'd765: data <= 32'hfd842783;
         'd766: data <= 32'h0047a703;         'd767: data <= 32'hfdc42783;
         'd768: data <= 32'h00e7a223;         'd769: data <= 32'hfd842783;
         'd770: data <= 32'hfec42703;         'd771: data <= 32'h00e7a223;
         'd772: data <= 32'hfd842783;         'd773: data <= 32'h0007a703;
         'd774: data <= 32'hfdc42783;         'd775: data <= 32'h00e7a023;
         'd776: data <= 32'hfd842783;         'd777: data <= 32'hfdc42703;
         'd778: data <= 32'h00e7a023;         'd779: data <= 32'hfdc42783;
         'd780: data <= 32'h00078513;         'd781: data <= 32'h02c12403;
         'd782: data <= 32'h03010113;         'd783: data <= 32'h00008067;
         'd784: data <= 32'hfe010113;         'd785: data <= 32'h00812e23;
         'd786: data <= 32'h02010413;         'd787: data <= 32'hfea42623;
         'd788: data <= 32'hfeb42423;         'd789: data <= 32'hfe842783;
         'd790: data <= 32'h00279783;         'd791: data <= 32'h0407c463;
         'd792: data <= 32'h0100006f;         'd793: data <= 32'hfec42783;
         'd794: data <= 32'h0007a783;         'd795: data <= 32'hfef42623;
         'd796: data <= 32'hfec42783;         'd797: data <= 32'h00078e63;
         'd798: data <= 32'hfec42783;         'd799: data <= 32'h0047a783;
         'd800: data <= 32'h00279703;         'd801: data <= 32'hfe842783;
         'd802: data <= 32'h00279783;         'd803: data <= 32'hfcf71ce3;
         'd804: data <= 32'hfec42783;         'd805: data <= 32'h0400006f;
         'd806: data <= 32'hfec42783;         'd807: data <= 32'h0007a783;
         'd808: data <= 32'hfef42623;         'd809: data <= 32'hfec42783;
         'd810: data <= 32'h02078463;         'd811: data <= 32'hfec42783;
         'd812: data <= 32'h0047a783;         'd813: data <= 32'h00079783;
         'd814: data <= 32'h01079793;         'd815: data <= 32'h0107d793;
         'd816: data <= 32'h0ff7f793;         'd817: data <= 32'hfe842703;
         'd818: data <= 32'h00071703;         'd819: data <= 32'hfce796e3;
         'd820: data <= 32'hfec42783;         'd821: data <= 32'h00078513;
         'd822: data <= 32'h01c12403;         'd823: data <= 32'h02010113;
         'd824: data <= 32'h00008067;         'd825: data <= 32'hfd010113;
         'd826: data <= 32'h02812623;         'd827: data <= 32'h03010413;
         'd828: data <= 32'hfca42e23;         'd829: data <= 32'hfe042623;
         'd830: data <= 32'h02c0006f;         'd831: data <= 32'hfdc42783;
         'd832: data <= 32'h0007a783;         'd833: data <= 32'hfef42423;
         'd834: data <= 32'hfdc42783;         'd835: data <= 32'hfec42703;
         'd836: data <= 32'h00e7a023;         'd837: data <= 32'hfdc42783;
         'd838: data <= 32'hfef42623;         'd839: data <= 32'hfe842783;
         'd840: data <= 32'hfcf42e23;         'd841: data <= 32'hfdc42783;
         'd842: data <= 32'hfc079ae3;         'd843: data <= 32'hfec42783;
         'd844: data <= 32'h00078513;         'd845: data <= 32'h02c12403;
         'd846: data <= 32'h03010113;         'd847: data <= 32'h00008067;
         'd848: data <= 32'hfb010113;         'd849: data <= 32'h04112623;
         'd850: data <= 32'h04812423;         'd851: data <= 32'h05010413;
         'd852: data <= 32'hfaa42e23;         'd853: data <= 32'hfab42c23;
         'd854: data <= 32'hfac42a23;         'd855: data <= 32'h00100793;
         'd856: data <= 32'hfcf42e23;         'd857: data <= 32'hfbc42783;
         'd858: data <= 32'hfef42623;         'd859: data <= 32'hfa042e23;
         'd860: data <= 32'hfe042023;         'd861: data <= 32'hfc042c23;
         'd862: data <= 32'h1880006f;         'd863: data <= 32'hfd842783;
         'd864: data <= 32'h00178793;         'd865: data <= 32'hfcf42c23;
         'd866: data <= 32'hfec42783;         'd867: data <= 32'hfef42423;
         'd868: data <= 32'hfc042a23;         'd869: data <= 32'hfc042623;
         'd870: data <= 32'h0300006f;         'd871: data <= 32'hfd442783;
         'd872: data <= 32'h00178793;         'd873: data <= 32'hfcf42a23;
         'd874: data <= 32'hfe842783;         'd875: data <= 32'h0007a783;
         'd876: data <= 32'hfef42423;         'd877: data <= 32'hfe842783;
         'd878: data <= 32'h02078063;         'd879: data <= 32'hfcc42783;
         'd880: data <= 32'h00178793;         'd881: data <= 32'hfcf42623;
         'd882: data <= 32'hfcc42703;         'd883: data <= 32'hfdc42783;
         'd884: data <= 32'hfcf746e3;         'd885: data <= 32'h0080006f;
         'd886: data <= 32'h00000013;         'd887: data <= 32'hfdc42783;
         'd888: data <= 32'hfcf42823;         'd889: data <= 32'h0fc0006f;
         'd890: data <= 32'hfd442783;         'd891: data <= 32'h02079463;
         'd892: data <= 32'hfe842783;         'd893: data <= 32'hfef42223;
         'd894: data <= 32'hfe842783;         'd895: data <= 32'h0007a783;
         'd896: data <= 32'hfef42423;         'd897: data <= 32'hfd042783;
         'd898: data <= 32'hfff78793;         'd899: data <= 32'hfcf42823;
         'd900: data <= 32'h0a80006f;         'd901: data <= 32'hfd042783;
         'd902: data <= 32'h00078663;         'd903: data <= 32'hfe842783;
         'd904: data <= 32'h02079463;         'd905: data <= 32'hfec42783;
         'd906: data <= 32'hfef42223;         'd907: data <= 32'hfec42783;
         'd908: data <= 32'h0007a783;         'd909: data <= 32'hfef42623;
         'd910: data <= 32'hfd442783;         'd911: data <= 32'hfff78793;
         'd912: data <= 32'hfcf42a23;         'd913: data <= 32'h0740006f;
         'd914: data <= 32'hfec42783;         'd915: data <= 32'h0047a703;
         'd916: data <= 32'hfe842783;         'd917: data <= 32'h0047a783;
         'd918: data <= 32'hfb842683;         'd919: data <= 32'hfb442603;
         'd920: data <= 32'h00078593;         'd921: data <= 32'h00070513;
         'd922: data <= 32'h000680e7;         'd923: data <= 32'h00050793;
         'd924: data <= 32'h02f04463;         'd925: data <= 32'hfec42783;
         'd926: data <= 32'hfef42223;         'd927: data <= 32'hfec42783;
         'd928: data <= 32'h0007a783;         'd929: data <= 32'hfef42623;
         'd930: data <= 32'hfd442783;         'd931: data <= 32'hfff78793;
         'd932: data <= 32'hfcf42a23;         'd933: data <= 32'h0240006f;
         'd934: data <= 32'hfe842783;         'd935: data <= 32'hfef42223;
         'd936: data <= 32'hfe842783;         'd937: data <= 32'h0007a783;
         'd938: data <= 32'hfef42423;         'd939: data <= 32'hfd042783;
         'd940: data <= 32'hfff78793;         'd941: data <= 32'hfcf42823;
         'd942: data <= 32'hfe042783;         'd943: data <= 32'h00078a63;
         'd944: data <= 32'hfe042783;         'd945: data <= 32'hfe442703;
         'd946: data <= 32'h00e7a023;         'd947: data <= 32'h00c0006f;
         'd948: data <= 32'hfe442783;         'd949: data <= 32'hfaf42e23;
         'd950: data <= 32'hfe442783;         'd951: data <= 32'hfef42023;
         'd952: data <= 32'hfd442783;         'd953: data <= 32'hf0f042e3;
         'd954: data <= 32'hfd042783;         'd955: data <= 32'h00f05663;
         'd956: data <= 32'hfe842783;         'd957: data <= 32'hee079ae3;
         'd958: data <= 32'hfe842783;         'd959: data <= 32'hfef42623;
         'd960: data <= 32'hfec42783;         'd961: data <= 32'he6079ce3;
         'd962: data <= 32'hfe042783;         'd963: data <= 32'h0007a023;
         'd964: data <= 32'hfd842703;         'd965: data <= 32'h00100793;
         'd966: data <= 32'h00e7c663;         'd967: data <= 32'hfbc42783;
         'd968: data <= 32'h0140006f;         'd969: data <= 32'hfdc42783;
         'd970: data <= 32'h00179793;         'd971: data <= 32'hfcf42e23;
         'd972: data <= 32'he35ff06f;         'd973: data <= 32'h00078513;
         'd974: data <= 32'h04c12083;         'd975: data <= 32'h04812403;
         'd976: data <= 32'h05010113;         'd977: data <= 32'h00008067;
         'd978: data <= 32'hfd010113;         'd979: data <= 32'h02112623;
         'd980: data <= 32'h02812423;         'd981: data <= 32'h03010413;
         'd982: data <= 32'hfca42e23;         'd983: data <= 32'hfdc42783;
         'd984: data <= 32'hfef42423;         'd985: data <= 32'hfe842783;
         'd986: data <= 32'h01c7a783;         'd987: data <= 32'hfef42223;
         'd988: data <= 32'hfe842783;         'd989: data <= 32'h02079c23;
         'd990: data <= 32'hfe842783;         'd991: data <= 32'h02079d23;
         'd992: data <= 32'hfe842783;         'd993: data <= 32'h02079e23;
         'd994: data <= 32'hfe842783;         'd995: data <= 32'h02079f23;
         'd996: data <= 32'hfe042623;         'd997: data <= 32'h0a00006f;
         'd998: data <= 32'h00100593;         'd999: data <= 32'hfe842503;
         'd1000: data <= 32'hce8ff0ef;         'd1001: data <= 32'h00050793;
         'd1002: data <= 32'hfef41123;         'd1003: data <= 32'hfe842783;
         'd1004: data <= 32'h0387d703;         'd1005: data <= 32'hfe245783;
         'd1006: data <= 32'h00070593;         'd1007: data <= 32'h00078513;
         'd1008: data <= 32'h6ac020ef;         'd1009: data <= 32'h00050793;
         'd1010: data <= 32'h00078713;         'd1011: data <= 32'hfe842783;
         'd1012: data <= 32'h02e79c23;         'd1013: data <= 32'hfff00593;
         'd1014: data <= 32'hfe842503;         'd1015: data <= 32'hcacff0ef;
         'd1016: data <= 32'h00050793;         'd1017: data <= 32'hfef41123;
         'd1018: data <= 32'hfe842783;         'd1019: data <= 32'h0387d703;
         'd1020: data <= 32'hfe245783;         'd1021: data <= 32'h00070593;
         'd1022: data <= 32'h00078513;         'd1023: data <= 32'h670020ef;
         'd1024: data <= 32'h00050793;         'd1025: data <= 32'h00078713;
         'd1026: data <= 32'hfe842783;         'd1027: data <= 32'h02e79c23;
         'd1028: data <= 32'hfec42783;         'd1029: data <= 32'h00079a63;
         'd1030: data <= 32'hfe842783;         'd1031: data <= 32'h0387d703;
         'd1032: data <= 32'hfe842783;         'd1033: data <= 32'h02e79d23;
         'd1034: data <= 32'hfec42783;         'd1035: data <= 32'h00178793;
         'd1036: data <= 32'hfef42623;         'd1037: data <= 32'hfec42703;
         'd1038: data <= 32'hfe442783;         'd1039: data <= 32'hf4f76ee3;
         'd1040: data <= 32'h00000793;         'd1041: data <= 32'h00078513;
         'd1042: data <= 32'h02c12083;         'd1043: data <= 32'h02812403;
         'd1044: data <= 32'h03010113;         'd1045: data <= 32'h00008067;
         'd1046: data <= 32'h81010113;         'd1047: data <= 32'h7e112623;
         'd1048: data <= 32'h7e812423;         'd1049: data <= 32'h7e912223;
         'd1050: data <= 32'h7f010413;         'd1051: data <= 32'hfa010113;
         'd1052: data <= 32'hfc042623;         'd1053: data <= 32'hfe041623;
         'd1054: data <= 32'hfe041523;         'd1055: data <= 32'hfff00793;
         'd1056: data <= 32'hfef41423;         'd1057: data <= 32'hfe041323;
         'd1058: data <= 32'hfc041b23;         'd1059: data <= 32'hfc840693;
         'd1060: data <= 32'hfcc40713;         'd1061: data <= 32'hf8440793;
         'd1062: data <= 32'h04278793;         'd1063: data <= 32'h00068613;
         'd1064: data <= 32'h00070593;         'd1065: data <= 32'h00078513;
         'd1066: data <= 32'h5fd030ef;         'd1067: data <= 32'h00100513;
         'd1068: data <= 32'h42c020ef;         'd1069: data <= 32'h00050793;
         'd1070: data <= 32'h01079793;         'd1071: data <= 32'h4107d793;
         'd1072: data <= 32'hf8f41223;         'd1073: data <= 32'h00200513;
         'd1074: data <= 32'h414020ef;         'd1075: data <= 32'h00050793;
         'd1076: data <= 32'h01079793;         'd1077: data <= 32'h4107d793;
         'd1078: data <= 32'hf8f41323;         'd1079: data <= 32'h00300513;
         'd1080: data <= 32'h3fc020ef;         'd1081: data <= 32'h00050793;
         'd1082: data <= 32'h01079793;         'd1083: data <= 32'h4107d793;
         'd1084: data <= 32'hf8f41423;         'd1085: data <= 32'h00400513;
         'd1086: data <= 32'h3e4020ef;         'd1087: data <= 32'h00050793;
         'd1088: data <= 32'hfaf42023;         'd1089: data <= 32'h00500513;
         'd1090: data <= 32'h3d4020ef;         'd1091: data <= 32'h00050793;
         'd1092: data <= 32'hfaf42223;         'd1093: data <= 32'hfa442783;
         'd1094: data <= 32'h00079663;         'd1095: data <= 32'h00700793;
         'd1096: data <= 32'hfaf42223;         'd1097: data <= 32'hf8441783;
         'd1098: data <= 32'h02079263;         'd1099: data <= 32'hf8641783;
         'd1100: data <= 32'h00079e63;         'd1101: data <= 32'hf8841783;
         'd1102: data <= 32'h00079a63;         'd1103: data <= 32'hf8041223;
         'd1104: data <= 32'hf8041323;         'd1105: data <= 32'h06600793;
         'd1106: data <= 32'hf8f41423;         'd1107: data <= 32'hf8441703;
         'd1108: data <= 32'h00100793;         'd1109: data <= 32'h02f71a63;
         'd1110: data <= 32'hf8641783;         'd1111: data <= 32'h02079663;
         'd1112: data <= 32'hf8841783;         'd1113: data <= 32'h02079263;
         'd1114: data <= 32'h000037b7;         'd1115: data <= 32'h41578793;
         'd1116: data <= 32'hf8f41223;         'd1117: data <= 32'h000037b7;
         'd1118: data <= 32'h41578793;         'd1119: data <= 32'hf8f41323;
         'd1120: data <= 32'h06600793;         'd1121: data <= 32'hf8f41423;
         'd1122: data <= 32'hfe041723;         'd1123: data <= 32'h1380006f;
         'd1124: data <= 32'hfee45703;         'd1125: data <= 32'h00070793;
         'd1126: data <= 32'h00579793;         'd1127: data <= 32'h40e787b3;
         'd1128: data <= 32'h00279793;         'd1129: data <= 32'h00e787b3;
         'd1130: data <= 32'h00479793;         'd1131: data <= 32'h00078693;
         'd1132: data <= 32'hfee45703;         'd1133: data <= 32'hfffff7b7;
         'd1134: data <= 32'h7c478793;         'd1135: data <= 32'hff040613;
         'd1136: data <= 32'h00f607b3;         'd1137: data <= 32'h00d786b3;
         'd1138: data <= 32'h00070793;         'd1139: data <= 32'h00479793;
         'd1140: data <= 32'h00e787b3;         'd1141: data <= 32'h00279793;
         'd1142: data <= 32'hff040713;         'd1143: data <= 32'h00f707b3;
         'd1144: data <= 32'hf8d7ae23;         'd1145: data <= 32'hfee45703;
         'd1146: data <= 32'h00070793;         'd1147: data <= 32'h00479793;
         'd1148: data <= 32'h00e787b3;         'd1149: data <= 32'h00279793;
         'd1150: data <= 32'hff040713;         'd1151: data <= 32'h00f707b3;
         'd1152: data <= 32'h7d000713;         'd1153: data <= 32'hfae7a623;
         'd1154: data <= 32'hfee45703;         'd1155: data <= 32'hf8441683;
         'd1156: data <= 32'h00070793;         'd1157: data <= 32'h00479793;
         'd1158: data <= 32'h00e787b3;         'd1159: data <= 32'h00279793;
         'd1160: data <= 32'hff040713;         'd1161: data <= 32'h00f707b3;
         'd1162: data <= 32'hf8d79a23;         'd1163: data <= 32'hfee45703;
         'd1164: data <= 32'hf8641683;         'd1165: data <= 32'h00070793;
         'd1166: data <= 32'h00479793;         'd1167: data <= 32'h00e787b3;
         'd1168: data <= 32'h00279793;         'd1169: data <= 32'hff040713;
         'd1170: data <= 32'h00f707b3;         'd1171: data <= 32'hf8d79b23;
         'd1172: data <= 32'hfee45703;         'd1173: data <= 32'hf8841683;
         'd1174: data <= 32'h00070793;         'd1175: data <= 32'h00479793;
         'd1176: data <= 32'h00e787b3;         'd1177: data <= 32'h00279793;
         'd1178: data <= 32'hff040713;         'd1179: data <= 32'h00f707b3;
         'd1180: data <= 32'hf8d79c23;         'd1181: data <= 32'hfee45703;
         'd1182: data <= 32'h00070793;         'd1183: data <= 32'h00479793;
         'd1184: data <= 32'h00e787b3;         'd1185: data <= 32'h00279793;
         'd1186: data <= 32'hff040713;         'd1187: data <= 32'h00f707b3;
         'd1188: data <= 32'hfc079a23;         'd1189: data <= 32'hfee45703;
         'd1190: data <= 32'hfa442683;         'd1191: data <= 32'h00070793;
         'd1192: data <= 32'h00479793;         'd1193: data <= 32'h00e787b3;
         'd1194: data <= 32'h00279793;         'd1195: data <= 32'hff040713;
         'd1196: data <= 32'h00f707b3;         'd1197: data <= 32'hfad7aa23;
         'd1198: data <= 32'hfee45783;         'd1199: data <= 32'h00178793;
         'd1200: data <= 32'hfef41723;         'd1201: data <= 32'hfee45783;
         'd1202: data <= 32'hec0784e3;         'd1203: data <= 32'hfe041723;
         'd1204: data <= 32'h0380006f;         'd1205: data <= 32'hfee45783;
         'd1206: data <= 32'h00100713;         'd1207: data <= 32'h00f717b3;
         'd1208: data <= 32'h00078713;         'd1209: data <= 32'hfa442783;
         'd1210: data <= 32'h00f777b3;         'd1211: data <= 32'h00078863;
         'd1212: data <= 32'hfea45783;         'd1213: data <= 32'h00178793;
         'd1214: data <= 32'hfef41523;         'd1215: data <= 32'hfee45783;
         'd1216: data <= 32'h00178793;         'd1217: data <= 32'hfef41723;
         'd1218: data <= 32'hfee45703;         'd1219: data <= 32'h00200793;
         'd1220: data <= 32'hfce7f2e3;         'd1221: data <= 32'hfe041723;
         'd1222: data <= 32'h0680006f;         'd1223: data <= 32'hfee45703;
         'd1224: data <= 32'h00070793;         'd1225: data <= 32'h00479793;
         'd1226: data <= 32'h00e787b3;         'd1227: data <= 32'h00279793;
         'd1228: data <= 32'hff040713;         'd1229: data <= 32'h00f707b3;
         'd1230: data <= 32'hfac7a783;         'd1231: data <= 32'hfea45703;
         'd1232: data <= 32'hfee45483;         'd1233: data <= 32'h00070593;
         'd1234: data <= 32'h00078513;         'd1235: data <= 32'h40d030ef;
         'd1236: data <= 32'h00050793;         'd1237: data <= 32'h00078713;
         'd1238: data <= 32'h00048793;         'd1239: data <= 32'h00479793;
         'd1240: data <= 32'h009787b3;         'd1241: data <= 32'h00279793;
         'd1242: data <= 32'hff040693;         'd1243: data <= 32'h00f687b3;
         'd1244: data <= 32'hfae7a623;         'd1245: data <= 32'hfee45783;
         'd1246: data <= 32'h00178793;         'd1247: data <= 32'hfef41723;
         'd1248: data <= 32'hfee45783;         'd1249: data <= 32'hf8078ce3;
         'd1250: data <= 32'hfe041723;         'd1251: data <= 32'h0c00006f;
         'd1252: data <= 32'hfee45783;         'd1253: data <= 32'h00100713;
         'd1254: data <= 32'h00f717b3;         'd1255: data <= 32'h00078713;
         'd1256: data <= 32'hfa442783;         'd1257: data <= 32'h00f777b3;
         'd1258: data <= 32'h08078c63;         'd1259: data <= 32'hfe042023;
         'd1260: data <= 32'h07c0006f;         'd1261: data <= 32'hfe042703;
         'd1262: data <= 32'h00070793;         'd1263: data <= 32'h00479793;
         'd1264: data <= 32'h00e787b3;         'd1265: data <= 32'h00279793;
         'd1266: data <= 32'hff040713;         'd1267: data <= 32'h00f707b3;
         'd1268: data <= 32'hf9c7a483;         'd1269: data <= 32'hf9c42783;
         'd1270: data <= 32'hfec45703;         'd1271: data <= 32'h00070593;
         'd1272: data <= 32'h00078513;         'd1273: data <= 32'h349030ef;
         'd1274: data <= 32'h00050793;         'd1275: data <= 32'h00078713;
         'd1276: data <= 32'hfee45783;         'd1277: data <= 32'h00178613;
         'd1278: data <= 32'h00e486b3;         'd1279: data <= 32'hfe042703;
         'd1280: data <= 32'h00070793;         'd1281: data <= 32'h00479793;
         'd1282: data <= 32'h00e787b3;         'd1283: data <= 32'h00c787b3;
         'd1284: data <= 32'h00279793;         'd1285: data <= 32'hff040713;
         'd1286: data <= 32'h00f707b3;         'd1287: data <= 32'hf8d7ae23;
         'd1288: data <= 32'hfe042783;         'd1289: data <= 32'h00178793;
         'd1290: data <= 32'hfef42023;         'd1291: data <= 32'hfe042783;
         'd1292: data <= 32'hf80782e3;         'd1293: data <= 32'hfec45783;
         'd1294: data <= 32'h00178793;         'd1295: data <= 32'hfef41623;
         'd1296: data <= 32'hfee45783;         'd1297: data <= 32'h00178793;
         'd1298: data <= 32'hfef41723;         'd1299: data <= 32'hfee45703;
         'd1300: data <= 32'h00200793;         'd1301: data <= 32'hf2e7fee3;
         'd1302: data <= 32'hfe041723;         'd1303: data <= 32'h1e80006f;
         'd1304: data <= 32'hfee45703;         'd1305: data <= 32'h00070793;
         'd1306: data <= 32'h00479793;         'd1307: data <= 32'h00e787b3;
         'd1308: data <= 32'h00279793;         'd1309: data <= 32'hff040713;
         'd1310: data <= 32'h00f707b3;         'd1311: data <= 32'hfb47a783;
         'd1312: data <= 32'h0017f793;         'd1313: data <= 32'h06078c63;
         'd1314: data <= 32'hf9c42683;         'd1315: data <= 32'hfee45703;
         'd1316: data <= 32'h00070793;         'd1317: data <= 32'h00479793;
         'd1318: data <= 32'h00e787b3;         'd1319: data <= 32'h00279793;
         'd1320: data <= 32'hff040713;         'd1321: data <= 32'h00f707b3;
         'd1322: data <= 32'hfa07a583;         'd1323: data <= 32'hfee45703;
         'd1324: data <= 32'h00070793;         'd1325: data <= 32'h00479793;
         'd1326: data <= 32'h00e787b3;         'd1327: data <= 32'h00279793;
         'd1328: data <= 32'hff040713;         'd1329: data <= 32'h00f707b3;
         'd1330: data <= 32'hf9479783;         'd1331: data <= 32'hfee45483;
         'd1332: data <= 32'h00078613;         'd1333: data <= 32'h00068513;
         'd1334: data <= 32'had4ff0ef;         'd1335: data <= 32'h00050713;
         'd1336: data <= 32'h00048793;         'd1337: data <= 32'h00479793;
         'd1338: data <= 32'h009787b3;         'd1339: data <= 32'h00279793;
         'd1340: data <= 32'hff040693;         'd1341: data <= 32'h00f687b3;
         'd1342: data <= 32'hfae7ac23;         'd1343: data <= 32'hfee45703;
         'd1344: data <= 32'h00070793;         'd1345: data <= 32'h00479793;
         'd1346: data <= 32'h00e787b3;         'd1347: data <= 32'h00279793;
         'd1348: data <= 32'hff040713;         'd1349: data <= 32'h00f707b3;
         'd1350: data <= 32'hfb47a783;         'd1351: data <= 32'h0027f793;
         'd1352: data <= 32'h0a078063;         'd1353: data <= 32'hf9c42503;
         'd1354: data <= 32'hfee45703;         'd1355: data <= 32'h00070793;
         'd1356: data <= 32'h00479793;         'd1357: data <= 32'h00e787b3;
         'd1358: data <= 32'h00279793;         'd1359: data <= 32'hff040713;
         'd1360: data <= 32'h00f707b3;         'd1361: data <= 32'hfa47a583;
         'd1362: data <= 32'hfee45703;         'd1363: data <= 32'h00070793;
         'd1364: data <= 32'h00479793;         'd1365: data <= 32'h00e787b3;
         'd1366: data <= 32'h00279793;         'd1367: data <= 32'hff040713;
         'd1368: data <= 32'h00f707b3;         'd1369: data <= 32'hf9479783;
         'd1370: data <= 32'h00078693;         'd1371: data <= 32'hfee45703;
         'd1372: data <= 32'h00070793;         'd1373: data <= 32'h00479793;
         'd1374: data <= 32'h00e787b3;         'd1375: data <= 32'h00279793;
         'd1376: data <= 32'hff040713;         'd1377: data <= 32'h00f707b3;
         'd1378: data <= 32'hf9679783;         'd1379: data <= 32'h01079793;
         'd1380: data <= 32'h00f6e633;         'd1381: data <= 32'hfee45703;
         'd1382: data <= 32'hf8440693;         'd1383: data <= 32'h00070793;
         'd1384: data <= 32'h00479793;         'd1385: data <= 32'h00e787b3;
         'd1386: data <= 32'h00279793;         'd1387: data <= 32'h02078793;
         'd1388: data <= 32'h00f687b3;         'd1389: data <= 32'h00878793;
         'd1390: data <= 32'h00078693;         'd1391: data <= 32'h415000ef;
         'd1392: data <= 32'hfee45703;         'd1393: data <= 32'h00070793;
         'd1394: data <= 32'h00479793;         'd1395: data <= 32'h00e787b3;
         'd1396: data <= 32'h00279793;         'd1397: data <= 32'hff040713;
         'd1398: data <= 32'h00f707b3;         'd1399: data <= 32'hfb47a783;
         'd1400: data <= 32'h0047f793;         'd1401: data <= 32'h04078a63;
         'd1402: data <= 32'hf9c42683;         'd1403: data <= 32'hfee45703;
         'd1404: data <= 32'h00070793;         'd1405: data <= 32'h00479793;
         'd1406: data <= 32'h00e787b3;         'd1407: data <= 32'h00279793;
         'd1408: data <= 32'hff040713;         'd1409: data <= 32'h00f707b3;
         'd1410: data <= 32'hf9479583;         'd1411: data <= 32'hfee45703;
         'd1412: data <= 32'h00070793;         'd1413: data <= 32'h00479793;
         'd1414: data <= 32'h00e787b3;         'd1415: data <= 32'h00279793;
         'd1416: data <= 32'hff040713;         'd1417: data <= 32'h00f707b3;
         'd1418: data <= 32'hfa87a783;         'd1419: data <= 32'h00078613;
         'd1420: data <= 32'h00068513;         'd1421: data <= 32'h045010ef;
         'd1422: data <= 32'hfee45783;         'd1423: data <= 32'h00178793;
         'd1424: data <= 32'hfef41723;         'd1425: data <= 32'hfee45783;
         'd1426: data <= 32'he0078ce3;         'd1427: data <= 32'hfa042783;
         'd1428: data <= 32'h0a079063;         'd1429: data <= 32'hfc042e23;
         'd1430: data <= 32'h00100793;         'd1431: data <= 32'hfaf42023;
         'd1432: data <= 32'h0440006f;         'd1433: data <= 32'hfa042703;
         'd1434: data <= 32'h00070793;         'd1435: data <= 32'h00279793;
         'd1436: data <= 32'h00e787b3;         'd1437: data <= 32'h00179793;
         'd1438: data <= 32'hfaf42023;         'd1439: data <= 32'h750030ef;
         'd1440: data <= 32'hf8440793;         'd1441: data <= 32'h00078513;
         'd1442: data <= 32'h8c1ff0ef;         'd1443: data <= 32'h770030ef;
         'd1444: data <= 32'h79c030ef;         'd1445: data <= 32'h00050793;
         'd1446: data <= 32'h00078513;         'd1447: data <= 32'h7c0030ef;
         'd1448: data <= 32'hfca42e23;         'd1449: data <= 32'hfdc42783;
         'd1450: data <= 32'hfa078ee3;         'd1451: data <= 32'hfdc42783;
         'd1452: data <= 32'hfcf42c23;         'd1453: data <= 32'hfd842783;
         'd1454: data <= 32'h00079663;         'd1455: data <= 32'h00100793;
         'd1456: data <= 32'hfcf42c23;         'd1457: data <= 32'hfa042483;
         'd1458: data <= 32'hfd842583;         'd1459: data <= 32'h00a00513;
         'd1460: data <= 32'h089030ef;         'd1461: data <= 32'h00050793;
         'd1462: data <= 32'h00178793;         'd1463: data <= 32'h00078593;
         'd1464: data <= 32'h00048513;         'd1465: data <= 32'h049030ef;
         'd1466: data <= 32'h00050793;         'd1467: data <= 32'hfaf42023;
         'd1468: data <= 32'h6dc030ef;         'd1469: data <= 32'hf8440793;
         'd1470: data <= 32'h00078513;         'd1471: data <= 32'h84dff0ef;
         'd1472: data <= 32'h6fc030ef;         'd1473: data <= 32'h728030ef;
         'd1474: data <= 32'hfca42823;         'd1475: data <= 32'hf8441783;
         'd1476: data <= 32'hfd645703;         'd1477: data <= 32'h00070593;
         'd1478: data <= 32'h00078513;         'd1479: data <= 32'h058020ef;
         'd1480: data <= 32'h00050793;         'd1481: data <= 32'hfcf41b23;
         'd1482: data <= 32'hf8641783;         'd1483: data <= 32'hfd645703;
         'd1484: data <= 32'h00070593;         'd1485: data <= 32'h00078513;
         'd1486: data <= 32'h03c020ef;         'd1487: data <= 32'h00050793;
         'd1488: data <= 32'hfcf41b23;         'd1489: data <= 32'hf8841783;
         'd1490: data <= 32'hfd645703;         'd1491: data <= 32'h00070593;
         'd1492: data <= 32'h00078513;         'd1493: data <= 32'h020020ef;
         'd1494: data <= 32'h00050793;         'd1495: data <= 32'hfcf41b23;
         'd1496: data <= 32'hf9c42783;         'd1497: data <= 32'h01079793;
         'd1498: data <= 32'h4107d793;         'd1499: data <= 32'hfd645703;
         'd1500: data <= 32'h00070593;         'd1501: data <= 32'h00078513;
         'd1502: data <= 32'h7fd010ef;         'd1503: data <= 32'h00050793;
         'd1504: data <= 32'hfcf41b23;         'd1505: data <= 32'hfd645783;
         'd1506: data <= 32'h0000f737;         'd1507: data <= 32'h9f570713;
         'd1508: data <= 32'h0ae78063;         'd1509: data <= 32'h0000f737;
         'd1510: data <= 32'h9f570713;         'd1511: data <= 32'h0cf74263;
         'd1512: data <= 32'h00009737;         'd1513: data <= 32'ha0270713;
         'd1514: data <= 32'h04e78263;         'd1515: data <= 32'h00009737;
         'd1516: data <= 32'ha0270713;         'd1517: data <= 32'h0af74663;
         'd1518: data <= 32'h00008737;         'd1519: data <= 32'hb0570713;
         'd1520: data <= 32'h04e78063;         'd1521: data <= 32'h00008737;
         'd1522: data <= 32'hb0570713;         'd1523: data <= 32'h08f74a63;
         'd1524: data <= 32'h00002737;         'd1525: data <= 32'h8f270713;
         'd1526: data <= 32'h06e78863;         'd1527: data <= 32'h00005737;
         'd1528: data <= 32'heaf70713;         'd1529: data <= 32'h02e78a63;
         'd1530: data <= 32'h0780006f;         'd1531: data <= 32'hfe041423;
         'd1532: data <= 32'h800057b7;         'd1533: data <= 32'h01c78513;
         'd1534: data <= 32'h2a8030ef;         'd1535: data <= 32'h0700006f;
         'd1536: data <= 32'h00100793;         'd1537: data <= 32'hfef41423;
         'd1538: data <= 32'h800057b7;         'd1539: data <= 32'h04c78513;
         'd1540: data <= 32'h290030ef;         'd1541: data <= 32'h0580006f;
         'd1542: data <= 32'h00200793;         'd1543: data <= 32'hfef41423;
         'd1544: data <= 32'h800057b7;         'd1545: data <= 32'h07878513;
         'd1546: data <= 32'h278030ef;         'd1547: data <= 32'h0400006f;
         'd1548: data <= 32'h00300793;         'd1549: data <= 32'hfef41423;
         'd1550: data <= 32'h800057b7;         'd1551: data <= 32'h0ac78513;
         'd1552: data <= 32'h260030ef;         'd1553: data <= 32'h0280006f;
         'd1554: data <= 32'h00400793;         'd1555: data <= 32'hfef41423;
         'd1556: data <= 32'h800057b7;         'd1557: data <= 32'h0dc78513;
         'd1558: data <= 32'h248030ef;         'd1559: data <= 32'h0100006f;
         'd1560: data <= 32'hfff00793;         'd1561: data <= 32'hfef41323;
         'd1562: data <= 32'h00000013;         'd1563: data <= 32'hfe841783;
         'd1564: data <= 32'h3807ce63;         'd1565: data <= 32'hfe041723;
         'd1566: data <= 32'h3880006f;         'd1567: data <= 32'hfee45703;
         'd1568: data <= 32'h00070793;         'd1569: data <= 32'h00479793;
         'd1570: data <= 32'h00e787b3;         'd1571: data <= 32'h00279793;
         'd1572: data <= 32'hff040713;         'd1573: data <= 32'h00f707b3;
         'd1574: data <= 32'hfc079a23;         'd1575: data <= 32'hfee45703;
         'd1576: data <= 32'h00070793;         'd1577: data <= 32'h00479793;
         'd1578: data <= 32'h00e787b3;         'd1579: data <= 32'h00279793;
         'd1580: data <= 32'hff040713;         'd1581: data <= 32'h00f707b3;
         'd1582: data <= 32'hfb47a783;         'd1583: data <= 32'h0017f793;
         'd1584: data <= 32'h0e078463;         'd1585: data <= 32'hfee45703;
         'd1586: data <= 32'h00070793;         'd1587: data <= 32'h00479793;
         'd1588: data <= 32'h00e787b3;         'd1589: data <= 32'h00279793;
         'd1590: data <= 32'hff040713;         'd1591: data <= 32'h00f707b3;
         'd1592: data <= 32'hfce7d703;         'd1593: data <= 32'hfe841783;
         'd1594: data <= 32'h100006b7;         'd1595: data <= 32'h00068693;
         'd1596: data <= 32'h00179793;         'd1597: data <= 32'h00f687b3;
         'd1598: data <= 32'h0007d783;         'd1599: data <= 32'h0af70663;
         'd1600: data <= 32'hfee45583;         'd1601: data <= 32'hfee45703;
         'd1602: data <= 32'h00070793;         'd1603: data <= 32'h00479793;
         'd1604: data <= 32'h00e787b3;         'd1605: data <= 32'h00279793;
         'd1606: data <= 32'hff040713;         'd1607: data <= 32'h00f707b3;
         'd1608: data <= 32'hfce7d783;         'd1609: data <= 32'h00078613;
         'd1610: data <= 32'hfe841783;         'd1611: data <= 32'h10000737;
         'd1612: data <= 32'h00070713;         'd1613: data <= 32'h00179793;
         'd1614: data <= 32'h00f707b3;         'd1615: data <= 32'h0007d783;
         'd1616: data <= 32'h00078693;         'd1617: data <= 32'h800057b7;
         'd1618: data <= 32'h10878513;         'd1619: data <= 32'h154030ef;
         'd1620: data <= 32'hfee45703;         'd1621: data <= 32'h00070793;
         'd1622: data <= 32'h00479793;         'd1623: data <= 32'h00e787b3;
         'd1624: data <= 32'h00279793;         'd1625: data <= 32'hff040693;
         'd1626: data <= 32'h00f687b3;         'd1627: data <= 32'hfd479783;
         'd1628: data <= 32'h01079793;         'd1629: data <= 32'h0107d793;
         'd1630: data <= 32'h00178793;         'd1631: data <= 32'h01079793;
         'd1632: data <= 32'h0107d793;         'd1633: data <= 32'h01079693;
         'd1634: data <= 32'h4106d693;         'd1635: data <= 32'h00070793;
         'd1636: data <= 32'h00479793;         'd1637: data <= 32'h00e787b3;
         'd1638: data <= 32'h00279793;         'd1639: data <= 32'hff040713;
         'd1640: data <= 32'h00f707b3;         'd1641: data <= 32'hfcd79a23;
         'd1642: data <= 32'hfee45703;         'd1643: data <= 32'h00070793;
         'd1644: data <= 32'h00479793;         'd1645: data <= 32'h00e787b3;
         'd1646: data <= 32'h00279793;         'd1647: data <= 32'hff040713;
         'd1648: data <= 32'h00f707b3;         'd1649: data <= 32'hfb47a783;
         'd1650: data <= 32'h0027f793;         'd1651: data <= 32'h0e078463;
         'd1652: data <= 32'hfee45703;         'd1653: data <= 32'h00070793;
         'd1654: data <= 32'h00479793;         'd1655: data <= 32'h00e787b3;
         'd1656: data <= 32'h00279793;         'd1657: data <= 32'hff040713;
         'd1658: data <= 32'h00f707b3;         'd1659: data <= 32'hfd07d703;
         'd1660: data <= 32'hfe841783;         'd1661: data <= 32'h100006b7;
         'd1662: data <= 32'h00c68693;         'd1663: data <= 32'h00179793;
         'd1664: data <= 32'h00f687b3;         'd1665: data <= 32'h0007d783;
         'd1666: data <= 32'h0af70663;         'd1667: data <= 32'hfee45583;
         'd1668: data <= 32'hfee45703;         'd1669: data <= 32'h00070793;
         'd1670: data <= 32'h00479793;         'd1671: data <= 32'h00e787b3;
         'd1672: data <= 32'h00279793;         'd1673: data <= 32'hff040713;
         'd1674: data <= 32'h00f707b3;         'd1675: data <= 32'hfd07d783;
         'd1676: data <= 32'h00078613;         'd1677: data <= 32'hfe841783;
         'd1678: data <= 32'h10000737;         'd1679: data <= 32'h00c70713;
         'd1680: data <= 32'h00179793;         'd1681: data <= 32'h00f707b3;
         'd1682: data <= 32'h0007d783;         'd1683: data <= 32'h00078693;
         'd1684: data <= 32'h800057b7;         'd1685: data <= 32'h13878513;
         'd1686: data <= 32'h048030ef;         'd1687: data <= 32'hfee45703;
         'd1688: data <= 32'h00070793;         'd1689: data <= 32'h00479793;
         'd1690: data <= 32'h00e787b3;         'd1691: data <= 32'h00279793;
         'd1692: data <= 32'hff040693;         'd1693: data <= 32'h00f687b3;
         'd1694: data <= 32'hfd479783;         'd1695: data <= 32'h01079793;
         'd1696: data <= 32'h0107d793;         'd1697: data <= 32'h00178793;
         'd1698: data <= 32'h01079793;         'd1699: data <= 32'h0107d793;
         'd1700: data <= 32'h01079693;         'd1701: data <= 32'h4106d693;
         'd1702: data <= 32'h00070793;         'd1703: data <= 32'h00479793;
         'd1704: data <= 32'h00e787b3;         'd1705: data <= 32'h00279793;
         'd1706: data <= 32'hff040713;         'd1707: data <= 32'h00f707b3;
         'd1708: data <= 32'hfcd79a23;         'd1709: data <= 32'hfee45703;
         'd1710: data <= 32'h00070793;         'd1711: data <= 32'h00479793;
         'd1712: data <= 32'h00e787b3;         'd1713: data <= 32'h00279793;
         'd1714: data <= 32'hff040713;         'd1715: data <= 32'h00f707b3;
         'd1716: data <= 32'hfb47a783;         'd1717: data <= 32'h0047f793;
         'd1718: data <= 32'h0e078063;         'd1719: data <= 32'hfee45703;
         'd1720: data <= 32'h00070793;         'd1721: data <= 32'h00479793;
         'd1722: data <= 32'h00e787b3;         'd1723: data <= 32'h00279793;
         'd1724: data <= 32'hff040713;         'd1725: data <= 32'h00f707b3;
         'd1726: data <= 32'hfd27d703;         'd1727: data <= 32'hfe841783;
         'd1728: data <= 32'h81818693;         'd1729: data <= 32'h00179793;
         'd1730: data <= 32'h00f687b3;         'd1731: data <= 32'h0007d783;
         'd1732: data <= 32'h0af70463;         'd1733: data <= 32'hfee45583;
         'd1734: data <= 32'hfee45703;         'd1735: data <= 32'h00070793;
         'd1736: data <= 32'h00479793;         'd1737: data <= 32'h00e787b3;
         'd1738: data <= 32'h00279793;         'd1739: data <= 32'hff040713;
         'd1740: data <= 32'h00f707b3;         'd1741: data <= 32'hfd27d783;
         'd1742: data <= 32'h00078613;         'd1743: data <= 32'hfe841783;
         'd1744: data <= 32'h81818713;         'd1745: data <= 32'h00179793;
         'd1746: data <= 32'h00f707b3;         'd1747: data <= 32'h0007d783;
         'd1748: data <= 32'h00078693;         'd1749: data <= 32'h800057b7;
         'd1750: data <= 32'h16c78513;         'd1751: data <= 32'h745020ef;
         'd1752: data <= 32'hfee45703;         'd1753: data <= 32'h00070793;
         'd1754: data <= 32'h00479793;         'd1755: data <= 32'h00e787b3;
         'd1756: data <= 32'h00279793;         'd1757: data <= 32'hff040693;
         'd1758: data <= 32'h00f687b3;         'd1759: data <= 32'hfd479783;
         'd1760: data <= 32'h01079793;         'd1761: data <= 32'h0107d793;
         'd1762: data <= 32'h00178793;         'd1763: data <= 32'h01079793;
         'd1764: data <= 32'h0107d793;         'd1765: data <= 32'h01079693;
         'd1766: data <= 32'h4106d693;         'd1767: data <= 32'h00070793;
         'd1768: data <= 32'h00479793;         'd1769: data <= 32'h00e787b3;
         'd1770: data <= 32'h00279793;         'd1771: data <= 32'hff040713;
         'd1772: data <= 32'h00f707b3;         'd1773: data <= 32'hfcd79a23;
         'd1774: data <= 32'hfee45703;         'd1775: data <= 32'h00070793;
         'd1776: data <= 32'h00479793;         'd1777: data <= 32'h00e787b3;
         'd1778: data <= 32'h00279793;         'd1779: data <= 32'hff040713;
         'd1780: data <= 32'h00f707b3;         'd1781: data <= 32'hfd479783;
         'd1782: data <= 32'h01079713;         'd1783: data <= 32'h01075713;
         'd1784: data <= 32'hfe645783;         'd1785: data <= 32'h00f707b3;
         'd1786: data <= 32'h01079793;         'd1787: data <= 32'h0107d793;
         'd1788: data <= 32'hfef41323;         'd1789: data <= 32'hfee45783;
         'd1790: data <= 32'h00178793;         'd1791: data <= 32'hfef41723;
         'd1792: data <= 32'hfee45703;         'd1793: data <= 32'h8741a783;
         'd1794: data <= 32'hc6f76ae3;         'd1795: data <= 32'h3b9010ef;
         'd1796: data <= 32'h00050793;         'd1797: data <= 32'h01079713;
         'd1798: data <= 32'h01075713;         'd1799: data <= 32'hfe645783;
         'd1800: data <= 32'h00f707b3;         'd1801: data <= 32'h01079793;
         'd1802: data <= 32'h0107d793;         'd1803: data <= 32'hfef41323;
         'd1804: data <= 32'hf9c42783;         'd1805: data <= 32'h00078593;
         'd1806: data <= 32'h800057b7;         'd1807: data <= 32'h19c78513;
         'd1808: data <= 32'h661020ef;         'd1809: data <= 32'hfd042583;
         'd1810: data <= 32'h800057b7;         'd1811: data <= 32'h1b478513;
         'd1812: data <= 32'h651020ef;         'd1813: data <= 32'hfd042503;
         'd1814: data <= 32'h204030ef;         'd1815: data <= 32'h00050793;
         'd1816: data <= 32'h00078593;         'd1817: data <= 32'h800057b7;
         'd1818: data <= 32'h1cc78513;         'd1819: data <= 32'h635020ef;
         'd1820: data <= 32'hfd042503;         'd1821: data <= 32'h1e8030ef;
         'd1822: data <= 32'h00050793;         'd1823: data <= 32'h04078663;
         'd1824: data <= 32'hfa042703;         'd1825: data <= 32'h8741a783;
         'd1826: data <= 32'h00078593;         'd1827: data <= 32'h00070513;
         'd1828: data <= 32'h29c030ef;         'd1829: data <= 32'h00050793;
         'd1830: data <= 32'h00078493;         'd1831: data <= 32'hfd042503;
         'd1832: data <= 32'h1bc030ef;         'd1833: data <= 32'h00050793;
         'd1834: data <= 32'h00078593;         'd1835: data <= 32'h00048513;
         'd1836: data <= 32'h2a8030ef;         'd1837: data <= 32'h00050793;
         'd1838: data <= 32'h00078593;         'd1839: data <= 32'h800057b7;
         'd1840: data <= 32'h1e478513;         'd1841: data <= 32'h5dd020ef;
         'd1842: data <= 32'hfd042503;         'd1843: data <= 32'h190030ef;
         'd1844: data <= 32'h00050713;         'd1845: data <= 32'h00900793;
         'd1846: data <= 32'h02e7e663;         'd1847: data <= 32'h800057b7;
         'd1848: data <= 32'h1fc78513;         'd1849: data <= 32'h5bd020ef;
         'd1850: data <= 32'hfe641783;         'd1851: data <= 32'h01079793;
         'd1852: data <= 32'h0107d793;         'd1853: data <= 32'h00178793;
         'd1854: data <= 32'h01079793;         'd1855: data <= 32'h0107d793;
         'd1856: data <= 32'hfef41323;         'd1857: data <= 32'hfa042703;
         'd1858: data <= 32'h8741a783;         'd1859: data <= 32'h00078593;
         'd1860: data <= 32'h00070513;         'd1861: data <= 32'h218030ef;
         'd1862: data <= 32'h00050793;         'd1863: data <= 32'h00078593;
         'd1864: data <= 32'h800057b7;         'd1865: data <= 32'h23c78513;
         'd1866: data <= 32'h579020ef;         'd1867: data <= 32'h800057b7;
         'd1868: data <= 32'h25478593;         'd1869: data <= 32'h800057b7;
         'd1870: data <= 32'h29878513;         'd1871: data <= 32'h565020ef;
         'd1872: data <= 32'h800057b7;         'd1873: data <= 32'h2b078593;
         'd1874: data <= 32'h800057b7;         'd1875: data <= 32'h39878513;
         'd1876: data <= 32'h551020ef;         'd1877: data <= 32'h800057b7;
         'd1878: data <= 32'h3b078593;         'd1879: data <= 32'h800057b7;
         'd1880: data <= 32'h3b878513;         'd1881: data <= 32'h53d020ef;
         'd1882: data <= 32'hfd645783;         'd1883: data <= 32'h00078593;
         'd1884: data <= 32'h800057b7;         'd1885: data <= 32'h3d078513;
         'd1886: data <= 32'h529020ef;         'd1887: data <= 32'hfa442783;
         'd1888: data <= 32'h0017f793;         'd1889: data <= 32'h04078e63;
         'd1890: data <= 32'hfe041723;         'd1891: data <= 32'h0480006f;
         'd1892: data <= 32'hfee45683;         'd1893: data <= 32'hfee45703;
         'd1894: data <= 32'h00070793;         'd1895: data <= 32'h00479793;
         'd1896: data <= 32'h00e787b3;         'd1897: data <= 32'h00279793;
         'd1898: data <= 32'hff040713;         'd1899: data <= 32'h00f707b3;
         'd1900: data <= 32'hfce7d783;         'd1901: data <= 32'h00078613;
         'd1902: data <= 32'h00068593;         'd1903: data <= 32'h800057b7;
         'd1904: data <= 32'h3ec78513;         'd1905: data <= 32'h4dd020ef;
         'd1906: data <= 32'hfee45783;         'd1907: data <= 32'h00178793;
         'd1908: data <= 32'hfef41723;         'd1909: data <= 32'hfee45703;
         'd1910: data <= 32'h8741a783;         'd1911: data <= 32'hfaf76ae3;
         'd1912: data <= 32'hfa442783;         'd1913: data <= 32'h0027f793;
         'd1914: data <= 32'h04078e63;         'd1915: data <= 32'hfe041723;
         'd1916: data <= 32'h0480006f;         'd1917: data <= 32'hfee45683;
         'd1918: data <= 32'hfee45703;         'd1919: data <= 32'h00070793;
         'd1920: data <= 32'h00479793;         'd1921: data <= 32'h00e787b3;
         'd1922: data <= 32'h00279793;         'd1923: data <= 32'hff040713;
         'd1924: data <= 32'h00f707b3;         'd1925: data <= 32'hfd07d783;
         'd1926: data <= 32'h00078613;         'd1927: data <= 32'h00068593;
         'd1928: data <= 32'h800057b7;         'd1929: data <= 32'h40878513;
         'd1930: data <= 32'h479020ef;         'd1931: data <= 32'hfee45783;
         'd1932: data <= 32'h00178793;         'd1933: data <= 32'hfef41723;
         'd1934: data <= 32'hfee45703;         'd1935: data <= 32'h8741a783;
         'd1936: data <= 32'hfaf76ae3;         'd1937: data <= 32'hfa442783;
         'd1938: data <= 32'h0047f793;         'd1939: data <= 32'h04078e63;
         'd1940: data <= 32'hfe041723;         'd1941: data <= 32'h0480006f;
         'd1942: data <= 32'hfee45683;         'd1943: data <= 32'hfee45703;
         'd1944: data <= 32'h00070793;         'd1945: data <= 32'h00479793;
         'd1946: data <= 32'h00e787b3;         'd1947: data <= 32'h00279793;
         'd1948: data <= 32'hff040713;         'd1949: data <= 32'h00f707b3;
         'd1950: data <= 32'hfd27d783;         'd1951: data <= 32'h00078613;
         'd1952: data <= 32'h00068593;         'd1953: data <= 32'h800057b7;
         'd1954: data <= 32'h42478513;         'd1955: data <= 32'h415020ef;
         'd1956: data <= 32'hfee45783;         'd1957: data <= 32'h00178793;
         'd1958: data <= 32'hfef41723;         'd1959: data <= 32'hfee45703;
         'd1960: data <= 32'h8741a783;         'd1961: data <= 32'hfaf76ae3;
         'd1962: data <= 32'hfe041723;         'd1963: data <= 32'h0480006f;
         'd1964: data <= 32'hfee45683;         'd1965: data <= 32'hfee45703;
         'd1966: data <= 32'h00070793;         'd1967: data <= 32'h00479793;
         'd1968: data <= 32'h00e787b3;         'd1969: data <= 32'h00279793;
         'd1970: data <= 32'hff040713;         'd1971: data <= 32'h00f707b3;
         'd1972: data <= 32'hfcc7d783;         'd1973: data <= 32'h00078613;
         'd1974: data <= 32'h00068593;         'd1975: data <= 32'h800057b7;
         'd1976: data <= 32'h44078513;         'd1977: data <= 32'h3bd020ef;
         'd1978: data <= 32'hfee45783;         'd1979: data <= 32'h00178793;
         'd1980: data <= 32'hfef41723;         'd1981: data <= 32'hfee45703;
         'd1982: data <= 32'h8741a783;         'd1983: data <= 32'hfaf76ae3;
         'd1984: data <= 32'hfe641783;         'd1985: data <= 32'h00079863;
         'd1986: data <= 32'h800057b7;         'd1987: data <= 32'h45c78513;
         'd1988: data <= 32'h391020ef;         'd1989: data <= 32'hfe641783;
         'd1990: data <= 32'h00f05863;         'd1991: data <= 32'h800057b7;
         'd1992: data <= 32'h4a878513;         'd1993: data <= 32'h37d020ef;
         'd1994: data <= 32'hfe641783;         'd1995: data <= 32'h0007d863;
         'd1996: data <= 32'h800057b7;         'd1997: data <= 32'h4bc78513;
         'd1998: data <= 32'h369020ef;         'd1999: data <= 32'hf8440793;
         'd2000: data <= 32'h04278793;         'd2001: data <= 32'h00078513;
         'd2002: data <= 32'h7c9020ef;         'd2003: data <= 32'h00000013;
         'd2004: data <= 32'h06010113;         'd2005: data <= 32'h7ec12083;
         'd2006: data <= 32'h7e812403;         'd2007: data <= 32'h7e412483;
         'd2008: data <= 32'h7f010113;         'd2009: data <= 32'h00008067;
         'd2010: data <= 32'hfc010113;         'd2011: data <= 32'h02112e23;
         'd2012: data <= 32'h02812c23;         'd2013: data <= 32'h04010413;
         'd2014: data <= 32'hfca42623;         'd2015: data <= 32'h00058793;
         'd2016: data <= 32'h00060713;         'd2017: data <= 32'hfcf41523;
         'd2018: data <= 32'h00070793;         'd2019: data <= 32'hfcf41423;
         'd2020: data <= 32'hfcc42783;         'd2021: data <= 32'h0007a783;
         'd2022: data <= 32'hfef42623;         'd2023: data <= 32'hfcc42783;
         'd2024: data <= 32'h00c7a783;         'd2025: data <= 32'hfef42423;
         'd2026: data <= 32'hfcc42783;         'd2027: data <= 32'h0047a783;
         'd2028: data <= 32'hfef42223;         'd2029: data <= 32'hfcc42783;
         'd2030: data <= 32'h0087a783;         'd2031: data <= 32'hfef42023;
         'd2032: data <= 32'hfca45783;         'd2033: data <= 32'hfcf41f23;
         'd2034: data <= 32'hfde41783;         'd2035: data <= 32'h00078713;
         'd2036: data <= 32'hfe042683;         'd2037: data <= 32'hfe442603;
         'd2038: data <= 32'hfe842583;         'd2039: data <= 32'hfec42503;
         'd2040: data <= 32'h03c000ef;         'd2041: data <= 32'h00050793;
         'd2042: data <= 32'h00078713;         'd2043: data <= 32'hfc845783;
         'd2044: data <= 32'h00078593;         'd2045: data <= 32'h00070513;
         'd2046: data <= 32'h77c010ef;         'd2047: data <= 32'h00050793;
         'd2048: data <= 32'hfcf41423;         'd2049: data <= 32'hfc845783;
         'd2050: data <= 32'h00078513;         'd2051: data <= 32'h03c12083;
         'd2052: data <= 32'h03812403;         'd2053: data <= 32'h04010113;
         'd2054: data <= 32'h00008067;         'd2055: data <= 32'hfc010113;
         'd2056: data <= 32'h02112e23;         'd2057: data <= 32'h02812c23;
         'd2058: data <= 32'h04010413;         'd2059: data <= 32'hfca42e23;
         'd2060: data <= 32'hfcb42c23;         'd2061: data <= 32'hfcc42a23;
         'd2062: data <= 32'hfcd42823;         'd2063: data <= 32'h00070793;
         'd2064: data <= 32'hfcf41723;         'd2065: data <= 32'hfe041723;
         'd2066: data <= 32'hfce45703;         'd2067: data <= 32'hfffff7b7;
         'd2068: data <= 32'h00f767b3;         'd2069: data <= 32'hfef41623;
         'd2070: data <= 32'hfce41783;         'd2071: data <= 32'h00078613;
         'd2072: data <= 32'hfd442583;         'd2073: data <= 32'hfdc42503;
         'd2074: data <= 32'h5ec000ef;         'd2075: data <= 32'hfce41783;
         'd2076: data <= 32'h00078693;         'd2077: data <= 32'hfd442603;
         'd2078: data <= 32'hfd842583;         'd2079: data <= 32'hfdc42503;
         'd2080: data <= 32'h4d0000ef;         'd2081: data <= 32'hfec41783;
         'd2082: data <= 32'h00078613;         'd2083: data <= 32'hfd842583;
         'd2084: data <= 32'hfdc42503;         'd2085: data <= 32'h398000ef;
         'd2086: data <= 32'h00050793;         'd2087: data <= 32'h00078713;
         'd2088: data <= 32'hfee45783;         'd2089: data <= 32'h00078593;
         'd2090: data <= 32'h00070513;         'd2091: data <= 32'h6c8010ef;
         'd2092: data <= 32'h00050793;         'd2093: data <= 32'hfef41723;
         'd2094: data <= 32'hfd042683;         'd2095: data <= 32'hfd442603;
         'd2096: data <= 32'hfd842583;         'd2097: data <= 32'hfdc42503;
         'd2098: data <= 32'h684000ef;         'd2099: data <= 32'hfec41783;
         'd2100: data <= 32'h00078613;         'd2101: data <= 32'hfd842583;
         'd2102: data <= 32'hfdc42503;         'd2103: data <= 32'h350000ef;
         'd2104: data <= 32'h00050793;         'd2105: data <= 32'h00078713;
         'd2106: data <= 32'hfee45783;         'd2107: data <= 32'h00078593;
         'd2108: data <= 32'h00070513;         'd2109: data <= 32'h680010ef;
         'd2110: data <= 32'h00050793;         'd2111: data <= 32'hfef41723;
         'd2112: data <= 32'hfd042683;         'd2113: data <= 32'hfd442603;
         'd2114: data <= 32'hfd842583;         'd2115: data <= 32'hfdc42503;
         'd2116: data <= 32'h754000ef;         'd2117: data <= 32'hfec41783;
         'd2118: data <= 32'h00078613;         'd2119: data <= 32'hfd842583;
         'd2120: data <= 32'hfdc42503;         'd2121: data <= 32'h308000ef;
         'd2122: data <= 32'h00050793;         'd2123: data <= 32'h00078713;
         'd2124: data <= 32'hfee45783;         'd2125: data <= 32'h00078593;
         'd2126: data <= 32'h00070513;         'd2127: data <= 32'h638010ef;
         'd2128: data <= 32'h00050793;         'd2129: data <= 32'hfef41723;
         'd2130: data <= 32'hfd042683;         'd2131: data <= 32'hfd442603;
         'd2132: data <= 32'hfd842583;         'd2133: data <= 32'hfdc42503;
         'd2134: data <= 32'h0ad000ef;         'd2135: data <= 32'hfec41783;
         'd2136: data <= 32'h00078613;         'd2137: data <= 32'hfd842583;
         'd2138: data <= 32'hfdc42503;         'd2139: data <= 32'h2c0000ef;
         'd2140: data <= 32'h00050793;         'd2141: data <= 32'h00078713;
         'd2142: data <= 32'hfee45783;         'd2143: data <= 32'h00078593;
         'd2144: data <= 32'h00070513;         'd2145: data <= 32'h5f0010ef;
         'd2146: data <= 32'h00050793;         'd2147: data <= 32'hfef41723;
         'd2148: data <= 32'hfce45783;         'd2149: data <= 32'h40f007b3;
         'd2150: data <= 32'h01079793;         'd2151: data <= 32'h0107d793;
         'd2152: data <= 32'h01079793;         'd2153: data <= 32'h4107d793;
         'd2154: data <= 32'h00078613;         'd2155: data <= 32'hfd442583;
         'd2156: data <= 32'hfdc42503;         'd2157: data <= 32'h4a0000ef;
         'd2158: data <= 32'hfee41783;         'd2159: data <= 32'h00078513;
         'd2160: data <= 32'h03c12083;         'd2161: data <= 32'h03812403;
         'd2162: data <= 32'h04010113;         'd2163: data <= 32'h00008067;
         'd2164: data <= 32'hfc010113;         'd2165: data <= 32'h02112e23;
         'd2166: data <= 32'h02812c23;         'd2167: data <= 32'h04010413;
         'd2168: data <= 32'hfca42623;         'd2169: data <= 32'hfcb42423;
         'd2170: data <= 32'hfcc42223;         'd2171: data <= 32'hfcd42023;
         'd2172: data <= 32'hfe042023;         'd2173: data <= 32'h00100793;
         'd2174: data <= 32'hfef42623;         'd2175: data <= 32'hfe042423;
         'd2176: data <= 32'hfe042223;         'd2177: data <= 32'hfc442783;
         'd2178: data <= 32'h02079a63;         'd2179: data <= 32'h00100793;
         'd2180: data <= 32'hfcf42223;         'd2181: data <= 32'h0280006f;
         'd2182: data <= 32'hfe842783;         'd2183: data <= 32'h00178793;
         'd2184: data <= 32'hfef42423;         'd2185: data <= 32'hfe842583;
         'd2186: data <= 32'hfe842503;         'd2187: data <= 32'h501020ef;
         'd2188: data <= 32'h00050793;         'd2189: data <= 32'h00379793;
         'd2190: data <= 32'hfef42223;         'd2191: data <= 32'hfe442703;
         'd2192: data <= 32'hfcc42783;         'd2193: data <= 32'hfcf76ae3;
         'd2194: data <= 32'hfe842783;         'd2195: data <= 32'hfff78793;
         'd2196: data <= 32'hfef42023;         'd2197: data <= 32'hfc842783;
         'd2198: data <= 32'hfff78793;         'd2199: data <= 32'hffc7f793;
         'd2200: data <= 32'h00478793;         'd2201: data <= 32'hfcf42e23;
         'd2202: data <= 32'hfe042583;         'd2203: data <= 32'hfe042503;
         'd2204: data <= 32'h4bd020ef;         'd2205: data <= 32'h00050793;
         'd2206: data <= 32'h00179793;         'd2207: data <= 32'hfdc42703;
         'd2208: data <= 32'h00f707b3;         'd2209: data <= 32'hfcf42c23;
         'd2210: data <= 32'hfe042423;         'd2211: data <= 32'h1240006f;
         'd2212: data <= 32'hfe042223;         'd2213: data <= 32'h1040006f;
         'd2214: data <= 32'hfc442583;         'd2215: data <= 32'hfec42503;
         'd2216: data <= 32'h48d020ef;         'd2217: data <= 32'h00050793;
         'd2218: data <= 32'h00078713;         'd2219: data <= 32'h41f75793;
         'd2220: data <= 32'h0107d793;         'd2221: data <= 32'h00f706b3;
         'd2222: data <= 32'h00010737;         'd2223: data <= 32'hfff70713;
         'd2224: data <= 32'h00e6f733;         'd2225: data <= 32'h40f707b3;
         'd2226: data <= 32'hfcf42223;         'd2227: data <= 32'hfc442783;
         'd2228: data <= 32'h01079713;         'd2229: data <= 32'h01075713;
         'd2230: data <= 32'hfec42783;         'd2231: data <= 32'h01079793;
         'd2232: data <= 32'h0107d793;         'd2233: data <= 32'h00f707b3;
         'd2234: data <= 32'h01079793;         'd2235: data <= 32'h0107d793;
         'd2236: data <= 32'hfcf41b23;         'd2237: data <= 32'hfe042583;
         'd2238: data <= 32'hfe842503;         'd2239: data <= 32'h431020ef;
         'd2240: data <= 32'h00050793;         'd2241: data <= 32'h00078713;
         'd2242: data <= 32'hfe442783;         'd2243: data <= 32'h00f707b3;
         'd2244: data <= 32'h00179793;         'd2245: data <= 32'hfd842703;
         'd2246: data <= 32'h00f707b3;         'd2247: data <= 32'hfd645703;
         'd2248: data <= 32'h00e79023;         'd2249: data <= 32'hfec42783;
         'd2250: data <= 32'h01079713;         'd2251: data <= 32'h01075713;
         'd2252: data <= 32'hfd645783;         'd2253: data <= 32'h00f707b3;
         'd2254: data <= 32'h01079793;         'd2255: data <= 32'h0107d793;
         'd2256: data <= 32'hfcf41b23;         'd2257: data <= 32'hfd645783;
         'd2258: data <= 32'h0ff7f793;         'd2259: data <= 32'hfcf41b23;
         'd2260: data <= 32'hfe042583;         'd2261: data <= 32'hfe842503;
         'd2262: data <= 32'h3d5020ef;         'd2263: data <= 32'h00050793;
         'd2264: data <= 32'h00078713;         'd2265: data <= 32'hfe442783;
         'd2266: data <= 32'h00f707b3;         'd2267: data <= 32'h00179793;
         'd2268: data <= 32'hfdc42703;         'd2269: data <= 32'h00f707b3;
         'd2270: data <= 32'hfd645703;         'd2271: data <= 32'h00e79023;
         'd2272: data <= 32'hfec42783;         'd2273: data <= 32'h00178793;
         'd2274: data <= 32'hfef42623;         'd2275: data <= 32'hfe442783;
         'd2276: data <= 32'h00178793;         'd2277: data <= 32'hfef42223;
         'd2278: data <= 32'hfe442703;         'd2279: data <= 32'hfe042783;
         'd2280: data <= 32'heef76ce3;         'd2281: data <= 32'hfe842783;
         'd2282: data <= 32'h00178793;         'd2283: data <= 32'hfef42423;
         'd2284: data <= 32'hfe842703;         'd2285: data <= 32'hfe042783;
         'd2286: data <= 32'hecf76ce3;         'd2287: data <= 32'hfc042783;
         'd2288: data <= 32'hfdc42703;         'd2289: data <= 32'h00e7a223;
         'd2290: data <= 32'hfc042783;         'd2291: data <= 32'hfd842703;
         'd2292: data <= 32'h00e7a423;         'd2293: data <= 32'hfe042583;
         'd2294: data <= 32'hfe042503;         'd2295: data <= 32'h351020ef;
         'd2296: data <= 32'h00050793;         'd2297: data <= 32'h00179793;
         'd2298: data <= 32'hfd842703;         'd2299: data <= 32'h00f707b3;
         'd2300: data <= 32'hfff78793;         'd2301: data <= 32'hffc7f793;
         'd2302: data <= 32'h00478793;         'd2303: data <= 32'h00078713;
         'd2304: data <= 32'hfc042783;         'd2305: data <= 32'h00e7a623;
         'd2306: data <= 32'hfe042703;         'd2307: data <= 32'hfc042783;
         'd2308: data <= 32'h00e7a023;         'd2309: data <= 32'hfe042783;
         'd2310: data <= 32'h00078513;         'd2311: data <= 32'h03c12083;
         'd2312: data <= 32'h03812403;         'd2313: data <= 32'h04010113;
         'd2314: data <= 32'h00008067;         'd2315: data <= 32'hfc010113;
         'd2316: data <= 32'h02112e23;         'd2317: data <= 32'h02812c23;
         'd2318: data <= 32'h04010413;         'd2319: data <= 32'hfca42623;
         'd2320: data <= 32'hfcb42423;         'd2321: data <= 32'h00060793;
         'd2322: data <= 32'hfcf41323;         'd2323: data <= 32'hfe042623;
         'd2324: data <= 32'hfe042423;         'd2325: data <= 32'hfc042c23;
         'd2326: data <= 32'hfe041323;         'd2327: data <= 32'hfe042023;
         'd2328: data <= 32'h0cc0006f;         'd2329: data <= 32'hfc042e23;
         'd2330: data <= 32'h0ac0006f;         'd2331: data <= 32'hfcc42583;
         'd2332: data <= 32'hfe042503;         'd2333: data <= 32'h2b9020ef;
         'd2334: data <= 32'h00050793;         'd2335: data <= 32'h00078713;
         'd2336: data <= 32'hfdc42783;         'd2337: data <= 32'h00f707b3;
         'd2338: data <= 32'h00279793;         'd2339: data <= 32'hfc842703;
         'd2340: data <= 32'h00f707b3;         'd2341: data <= 32'h0007a783;
         'd2342: data <= 32'hfcf42c23;         'd2343: data <= 32'hfec42703;
         'd2344: data <= 32'hfd842783;         'd2345: data <= 32'h00f707b3;
         'd2346: data <= 32'hfef42623;         'd2347: data <= 32'hfc641783;
         'd2348: data <= 32'hfec42703;         'd2349: data <= 32'h02e7d063;
         'd2350: data <= 32'hfe645783;         'd2351: data <= 32'h00a78793;
         'd2352: data <= 32'h01079793;         'd2353: data <= 32'h0107d793;
         'd2354: data <= 32'hfef41323;         'd2355: data <= 32'hfe042623;
         'd2356: data <= 32'h0300006f;         'd2357: data <= 32'hfd842703;
         'd2358: data <= 32'hfe842783;         'd2359: data <= 32'h00e7a7b3;
         'd2360: data <= 32'h0ff7f793;         'd2361: data <= 32'h01079713;
         'd2362: data <= 32'h01075713;         'd2363: data <= 32'hfe645783;
         'd2364: data <= 32'h00f707b3;         'd2365: data <= 32'h01079793;
         'd2366: data <= 32'h0107d793;         'd2367: data <= 32'hfef41323;
         'd2368: data <= 32'hfd842783;         'd2369: data <= 32'hfef42423;
         'd2370: data <= 32'hfdc42783;         'd2371: data <= 32'h00178793;
         'd2372: data <= 32'hfcf42e23;         'd2373: data <= 32'hfdc42703;
         'd2374: data <= 32'hfcc42783;         'd2375: data <= 32'hf4f768e3;
         'd2376: data <= 32'hfe042783;         'd2377: data <= 32'h00178793;
         'd2378: data <= 32'hfef42023;         'd2379: data <= 32'hfe042703;
         'd2380: data <= 32'hfcc42783;         'd2381: data <= 32'hf2f768e3;
         'd2382: data <= 32'hfe641783;         'd2383: data <= 32'h00078513;
         'd2384: data <= 32'h03c12083;         'd2385: data <= 32'h03812403;
         'd2386: data <= 32'h04010113;         'd2387: data <= 32'h00008067;
         'd2388: data <= 32'hfc010113;         'd2389: data <= 32'h02112e23;
         'd2390: data <= 32'h02812c23;         'd2391: data <= 32'h02912a23;
         'd2392: data <= 32'h03212823;         'd2393: data <= 32'h03312623;
         'd2394: data <= 32'h04010413;         'd2395: data <= 32'hfca42623;
         'd2396: data <= 32'hfcb42423;         'd2397: data <= 32'hfcc42223;
         'd2398: data <= 32'h00068793;         'd2399: data <= 32'hfcf41123;
         'd2400: data <= 32'hfc042e23;         'd2401: data <= 32'h0a00006f;
         'd2402: data <= 32'hfc042c23;         'd2403: data <= 32'h0800006f;
         'd2404: data <= 32'hfcc42583;         'd2405: data <= 32'hfdc42503;
         'd2406: data <= 32'h195020ef;         'd2407: data <= 32'h00050793;
         'd2408: data <= 32'h00078713;         'd2409: data <= 32'hfd842783;
         'd2410: data <= 32'h00f707b3;         'd2411: data <= 32'h00179793;
         'd2412: data <= 32'hfc442703;         'd2413: data <= 32'h00f707b3;
         'd2414: data <= 32'h00079783;         'd2415: data <= 32'h00078993;
         'd2416: data <= 32'hfc241903;         'd2417: data <= 32'hfcc42583;
         'd2418: data <= 32'hfdc42503;         'd2419: data <= 32'h161020ef;
         'd2420: data <= 32'h00050793;         'd2421: data <= 32'h00078713;
         'd2422: data <= 32'hfd842783;         'd2423: data <= 32'h00f707b3;
         'd2424: data <= 32'h00279793;         'd2425: data <= 32'hfc842703;
         'd2426: data <= 32'h00f704b3;         'd2427: data <= 32'h00090593;
         'd2428: data <= 32'h00098513;         'd2429: data <= 32'h139020ef;
         'd2430: data <= 32'h00050793;         'd2431: data <= 32'h00f4a023;
         'd2432: data <= 32'hfd842783;         'd2433: data <= 32'h00178793;
         'd2434: data <= 32'hfcf42c23;         'd2435: data <= 32'hfd842703;
         'd2436: data <= 32'hfcc42783;         'd2437: data <= 32'hf6f76ee3;
         'd2438: data <= 32'hfdc42783;         'd2439: data <= 32'h00178793;
         'd2440: data <= 32'hfcf42e23;         'd2441: data <= 32'hfdc42703;
         'd2442: data <= 32'hfcc42783;         'd2443: data <= 32'hf4f76ee3;
         'd2444: data <= 32'h00000013;         'd2445: data <= 32'h00000013;
         'd2446: data <= 32'h03c12083;         'd2447: data <= 32'h03812403;
         'd2448: data <= 32'h03412483;         'd2449: data <= 32'h03012903;
         'd2450: data <= 32'h02c12983;         'd2451: data <= 32'h04010113;
         'd2452: data <= 32'h00008067;         'd2453: data <= 32'hfd010113;
         'd2454: data <= 32'h02112623;         'd2455: data <= 32'h02812423;
         'd2456: data <= 32'h02912223;         'd2457: data <= 32'h03010413;
         'd2458: data <= 32'hfca42e23;         'd2459: data <= 32'hfcb42c23;
         'd2460: data <= 32'h00060793;         'd2461: data <= 32'hfcf41b23;
         'd2462: data <= 32'hfe042623;         'd2463: data <= 32'h0a80006f;
         'd2464: data <= 32'hfe042423;         'd2465: data <= 32'h0880006f;
         'd2466: data <= 32'hfdc42583;         'd2467: data <= 32'hfec42503;
         'd2468: data <= 32'h09d020ef;         'd2469: data <= 32'h00050793;
         'd2470: data <= 32'h00078713;         'd2471: data <= 32'hfe842783;
         'd2472: data <= 32'h00f707b3;         'd2473: data <= 32'h00179793;
         'd2474: data <= 32'hfd842703;         'd2475: data <= 32'h00f707b3;
         'd2476: data <= 32'h00079783;         'd2477: data <= 32'h01079713;
         'd2478: data <= 32'h01075713;         'd2479: data <= 32'hfd645783;
         'd2480: data <= 32'h00f707b3;         'd2481: data <= 32'h01079493;
         'd2482: data <= 32'h0104d493;         'd2483: data <= 32'hfdc42583;
         'd2484: data <= 32'hfec42503;         'd2485: data <= 32'h059020ef;
         'd2486: data <= 32'h00050793;         'd2487: data <= 32'h00078713;
         'd2488: data <= 32'hfe842783;         'd2489: data <= 32'h00f707b3;
         'd2490: data <= 32'h00179793;         'd2491: data <= 32'hfd842703;
         'd2492: data <= 32'h00f707b3;         'd2493: data <= 32'h01049713;
         'd2494: data <= 32'h41075713;         'd2495: data <= 32'h00e79023;
         'd2496: data <= 32'hfe842783;         'd2497: data <= 32'h00178793;
         'd2498: data <= 32'hfef42423;         'd2499: data <= 32'hfe842703;
         'd2500: data <= 32'hfdc42783;         'd2501: data <= 32'hf6f76ae3;
         'd2502: data <= 32'hfec42783;         'd2503: data <= 32'h00178793;
         'd2504: data <= 32'hfef42623;         'd2505: data <= 32'hfec42703;
         'd2506: data <= 32'hfdc42783;         'd2507: data <= 32'hf4f76ae3;
         'd2508: data <= 32'h00000013;         'd2509: data <= 32'h00000013;
         'd2510: data <= 32'h02c12083;         'd2511: data <= 32'h02812403;
         'd2512: data <= 32'h02412483;         'd2513: data <= 32'h03010113;
         'd2514: data <= 32'h00008067;         'd2515: data <= 32'hfd010113;
         'd2516: data <= 32'h02112623;         'd2517: data <= 32'h02812423;
         'd2518: data <= 32'h02912223;         'd2519: data <= 32'h03010413;
         'd2520: data <= 32'hfca42e23;         'd2521: data <= 32'hfcb42c23;
         'd2522: data <= 32'hfcc42a23;         'd2523: data <= 32'hfcd42823;
         'd2524: data <= 32'hfe042623;         'd2525: data <= 32'h0c80006f;
         'd2526: data <= 32'hfec42783;         'd2527: data <= 32'h00279793;
         'd2528: data <= 32'hfd842703;         'd2529: data <= 32'h00f707b3;
         'd2530: data <= 32'h0007a023;         'd2531: data <= 32'hfe042423;
         'd2532: data <= 32'h0940006f;         'd2533: data <= 32'hfec42783;
         'd2534: data <= 32'h00279793;         'd2535: data <= 32'hfd842703;
         'd2536: data <= 32'h00f707b3;         'd2537: data <= 32'h0007a483;
         'd2538: data <= 32'hfdc42583;         'd2539: data <= 32'hfec42503;
         'd2540: data <= 32'h77c020ef;         'd2541: data <= 32'h00050793;
         'd2542: data <= 32'h00078713;         'd2543: data <= 32'hfe842783;
         'd2544: data <= 32'h00f707b3;         'd2545: data <= 32'h00179793;
         'd2546: data <= 32'hfd442703;         'd2547: data <= 32'h00f707b3;
         'd2548: data <= 32'h00079783;         'd2549: data <= 32'h00078693;
         'd2550: data <= 32'hfe842783;         'd2551: data <= 32'h00179793;
         'd2552: data <= 32'hfd042703;         'd2553: data <= 32'h00f707b3;
         'd2554: data <= 32'h00079783;         'd2555: data <= 32'h00078593;
         'd2556: data <= 32'h00068513;         'd2557: data <= 32'h738020ef;
         'd2558: data <= 32'h00050793;         'd2559: data <= 32'h00078693;
         'd2560: data <= 32'hfec42783;         'd2561: data <= 32'h00279793;
         'd2562: data <= 32'hfd842703;         'd2563: data <= 32'h00f707b3;
         'd2564: data <= 32'h00d48733;         'd2565: data <= 32'h00e7a023;
         'd2566: data <= 32'hfe842783;         'd2567: data <= 32'h00178793;
         'd2568: data <= 32'hfef42423;         'd2569: data <= 32'hfe842703;
         'd2570: data <= 32'hfdc42783;         'd2571: data <= 32'hf6f764e3;
         'd2572: data <= 32'hfec42783;         'd2573: data <= 32'h00178793;
         'd2574: data <= 32'hfef42623;         'd2575: data <= 32'hfec42703;
         'd2576: data <= 32'hfdc42783;         'd2577: data <= 32'hf2f76ae3;
         'd2578: data <= 32'h00000013;         'd2579: data <= 32'h00000013;
         'd2580: data <= 32'h02c12083;         'd2581: data <= 32'h02812403;
         'd2582: data <= 32'h02412483;         'd2583: data <= 32'h03010113;
         'd2584: data <= 32'h00008067;         'd2585: data <= 32'hfd010113;
         'd2586: data <= 32'h02112623;         'd2587: data <= 32'h02812423;
         'd2588: data <= 32'h02912223;         'd2589: data <= 32'h03212023;
         'd2590: data <= 32'h03010413;         'd2591: data <= 32'hfca42e23;
         'd2592: data <= 32'hfcb42c23;         'd2593: data <= 32'hfcc42a23;
         'd2594: data <= 32'hfcd42823;         'd2595: data <= 32'hfe042623;
         'd2596: data <= 32'h1480006f;         'd2597: data <= 32'hfe042423;
         'd2598: data <= 32'h1280006f;         'd2599: data <= 32'hfdc42583;
         'd2600: data <= 32'hfec42503;         'd2601: data <= 32'h688020ef;
         'd2602: data <= 32'h00050793;         'd2603: data <= 32'h00078713;
         'd2604: data <= 32'hfe842783;         'd2605: data <= 32'h00f707b3;
         'd2606: data <= 32'h00279793;         'd2607: data <= 32'hfd842703;
         'd2608: data <= 32'h00f707b3;         'd2609: data <= 32'h0007a023;
         'd2610: data <= 32'hfe042223;         'd2611: data <= 32'h0dc0006f;
         'd2612: data <= 32'hfdc42583;         'd2613: data <= 32'hfec42503;
         'd2614: data <= 32'h654020ef;         'd2615: data <= 32'h00050793;
         'd2616: data <= 32'h00078713;         'd2617: data <= 32'hfe842783;
         'd2618: data <= 32'h00f707b3;         'd2619: data <= 32'h00279793;
         'd2620: data <= 32'hfd842703;         'd2621: data <= 32'h00f707b3;
         'd2622: data <= 32'h0007a483;         'd2623: data <= 32'hfdc42583;
         'd2624: data <= 32'hfec42503;         'd2625: data <= 32'h628020ef;
         'd2626: data <= 32'h00050793;         'd2627: data <= 32'h00078713;
         'd2628: data <= 32'hfe442783;         'd2629: data <= 32'h00f707b3;
         'd2630: data <= 32'h00179793;         'd2631: data <= 32'hfd442703;
         'd2632: data <= 32'h00f707b3;         'd2633: data <= 32'h00079783;
         'd2634: data <= 32'h00078913;         'd2635: data <= 32'hfdc42583;
         'd2636: data <= 32'hfe442503;         'd2637: data <= 32'h5f8020ef;
         'd2638: data <= 32'h00050793;         'd2639: data <= 32'h00078713;
         'd2640: data <= 32'hfe842783;         'd2641: data <= 32'h00f707b3;
         'd2642: data <= 32'h00179793;         'd2643: data <= 32'hfd042703;
         'd2644: data <= 32'h00f707b3;         'd2645: data <= 32'h00079783;
         'd2646: data <= 32'h00078593;         'd2647: data <= 32'h00090513;
         'd2648: data <= 32'h5cc020ef;         'd2649: data <= 32'h00050793;
         'd2650: data <= 32'h00078913;         'd2651: data <= 32'hfdc42583;
         'd2652: data <= 32'hfec42503;         'd2653: data <= 32'h5b8020ef;
         'd2654: data <= 32'h00050793;         'd2655: data <= 32'h00078713;
         'd2656: data <= 32'hfe842783;         'd2657: data <= 32'h00f707b3;
         'd2658: data <= 32'h00279793;         'd2659: data <= 32'hfd842703;
         'd2660: data <= 32'h00f707b3;         'd2661: data <= 32'h01248733;
         'd2662: data <= 32'h00e7a023;         'd2663: data <= 32'hfe442783;
         'd2664: data <= 32'h00178793;         'd2665: data <= 32'hfef42223;
         'd2666: data <= 32'hfe442703;         'd2667: data <= 32'hfdc42783;
         'd2668: data <= 32'hf2f760e3;         'd2669: data <= 32'hfe842783;
         'd2670: data <= 32'h00178793;         'd2671: data <= 32'hfef42423;
         'd2672: data <= 32'hfe842703;         'd2673: data <= 32'hfdc42783;
         'd2674: data <= 32'hecf76ae3;         'd2675: data <= 32'hfec42783;
         'd2676: data <= 32'h00178793;         'd2677: data <= 32'hfef42623;
         'd2678: data <= 32'hfec42703;         'd2679: data <= 32'hfdc42783;
         'd2680: data <= 32'heaf76ae3;         'd2681: data <= 32'h00000013;
         'd2682: data <= 32'h00000013;         'd2683: data <= 32'h02c12083;
         'd2684: data <= 32'h02812403;         'd2685: data <= 32'h02412483;
         'd2686: data <= 32'h02012903;         'd2687: data <= 32'h03010113;
         'd2688: data <= 32'h00008067;         'd2689: data <= 32'hfd010113;
         'd2690: data <= 32'h02112623;         'd2691: data <= 32'h02812423;
         'd2692: data <= 32'h02912223;         'd2693: data <= 32'h03010413;
         'd2694: data <= 32'hfca42e23;         'd2695: data <= 32'hfcb42c23;
         'd2696: data <= 32'hfcc42a23;         'd2697: data <= 32'hfcd42823;
         'd2698: data <= 32'hfe042623;         'd2699: data <= 32'h1780006f;
         'd2700: data <= 32'hfe042423;         'd2701: data <= 32'h1580006f;
         'd2702: data <= 32'hfdc42583;         'd2703: data <= 32'hfec42503;
         'd2704: data <= 32'h4ec020ef;         'd2705: data <= 32'h00050793;
         'd2706: data <= 32'h00078713;         'd2707: data <= 32'hfe842783;
         'd2708: data <= 32'h00f707b3;         'd2709: data <= 32'h00279793;
         'd2710: data <= 32'hfd842703;         'd2711: data <= 32'h00f707b3;
         'd2712: data <= 32'h0007a023;         'd2713: data <= 32'hfe042223;
         'd2714: data <= 32'h10c0006f;         'd2715: data <= 32'hfdc42583;
         'd2716: data <= 32'hfec42503;         'd2717: data <= 32'h4b8020ef;
         'd2718: data <= 32'h00050793;         'd2719: data <= 32'h00078713;
         'd2720: data <= 32'hfe442783;         'd2721: data <= 32'h00f707b3;
         'd2722: data <= 32'h00179793;         'd2723: data <= 32'hfd442703;
         'd2724: data <= 32'h00f707b3;         'd2725: data <= 32'h00079783;
         'd2726: data <= 32'h00078493;         'd2727: data <= 32'hfdc42583;
         'd2728: data <= 32'hfe442503;         'd2729: data <= 32'h488020ef;
         'd2730: data <= 32'h00050793;         'd2731: data <= 32'h00078713;
         'd2732: data <= 32'hfe842783;         'd2733: data <= 32'h00f707b3;
         'd2734: data <= 32'h00179793;         'd2735: data <= 32'hfd042703;
         'd2736: data <= 32'h00f707b3;         'd2737: data <= 32'h00079783;
         'd2738: data <= 32'h00078593;         'd2739: data <= 32'h00048513;
         'd2740: data <= 32'h45c020ef;         'd2741: data <= 32'h00050793;
         'd2742: data <= 32'hfef42023;         'd2743: data <= 32'hfdc42583;
         'd2744: data <= 32'hfec42503;         'd2745: data <= 32'h448020ef;
         'd2746: data <= 32'h00050793;         'd2747: data <= 32'h00078713;
         'd2748: data <= 32'hfe842783;         'd2749: data <= 32'h00f707b3;
         'd2750: data <= 32'h00279793;         'd2751: data <= 32'hfd842703;
         'd2752: data <= 32'h00f707b3;         'd2753: data <= 32'h0007a783;
         'd2754: data <= 32'h00078493;         'd2755: data <= 32'hfe042783;
         'd2756: data <= 32'h4027d793;         'd2757: data <= 32'h00f7f713;
         'd2758: data <= 32'hfe042783;         'd2759: data <= 32'h4057d793;
         'd2760: data <= 32'h07f7f793;         'd2761: data <= 32'h00078593;
         'd2762: data <= 32'h00070513;         'd2763: data <= 32'h400020ef;
         'd2764: data <= 32'h00050793;         'd2765: data <= 32'h00f484b3;
         'd2766: data <= 32'hfdc42583;         'd2767: data <= 32'hfec42503;
         'd2768: data <= 32'h3ec020ef;         'd2769: data <= 32'h00050793;
         'd2770: data <= 32'h00078713;         'd2771: data <= 32'hfe842783;
         'd2772: data <= 32'h00f707b3;         'd2773: data <= 32'h00279793;
         'd2774: data <= 32'hfd842703;         'd2775: data <= 32'h00f707b3;
         'd2776: data <= 32'h00048713;         'd2777: data <= 32'h00e7a023;
         'd2778: data <= 32'hfe442783;         'd2779: data <= 32'h00178793;
         'd2780: data <= 32'hfef42223;         'd2781: data <= 32'hfe442703;
         'd2782: data <= 32'hfdc42783;         'd2783: data <= 32'heef768e3;
         'd2784: data <= 32'hfe842783;         'd2785: data <= 32'h00178793;
         'd2786: data <= 32'hfef42423;         'd2787: data <= 32'hfe842703;
         'd2788: data <= 32'hfdc42783;         'd2789: data <= 32'heaf762e3;
         'd2790: data <= 32'hfec42783;         'd2791: data <= 32'h00178793;
         'd2792: data <= 32'hfef42623;         'd2793: data <= 32'hfec42703;
         'd2794: data <= 32'hfdc42783;         'd2795: data <= 32'he8f762e3;
         'd2796: data <= 32'h00000013;         'd2797: data <= 32'h00000013;
         'd2798: data <= 32'h02c12083;         'd2799: data <= 32'h02812403;
         'd2800: data <= 32'h02412483;         'd2801: data <= 32'h03010113;
         'd2802: data <= 32'h00008067;         'd2803: data <= 32'hf9010113;
         'd2804: data <= 32'h06112623;         'd2805: data <= 32'h06812423;
         'd2806: data <= 32'h07010413;         'd2807: data <= 32'hf8a42e23;
         'd2808: data <= 32'hf8b42c23;         'd2809: data <= 32'h00060593;
         'd2810: data <= 32'h00068613;         'd2811: data <= 32'h00070693;
         'd2812: data <= 32'h00078713;         'd2813: data <= 32'h00058793;
         'd2814: data <= 32'hf8f41b23;         'd2815: data <= 32'h00060793;
         'd2816: data <= 32'hf8f41a23;         'd2817: data <= 32'h00068793;
         'd2818: data <= 32'hf8f41923;         'd2819: data <= 32'h00070793;
         'd2820: data <= 32'hf8f41823;         'd2821: data <= 32'hf9842783;
         'd2822: data <= 32'hfaf42023;         'd2823: data <= 32'hfe042623;
         'd2824: data <= 32'h04c0006f;         'd2825: data <= 32'hfec42783;
         'd2826: data <= 32'h00279793;         'd2827: data <= 32'hff040713;
         'd2828: data <= 32'h00f707b3;         'd2829: data <= 32'hfa07aa23;
         'd2830: data <= 32'hfec42783;         'd2831: data <= 32'h00279793;
         'd2832: data <= 32'hff040713;         'd2833: data <= 32'h00f707b3;
         'd2834: data <= 32'hfb47a703;         'd2835: data <= 32'hfec42783;
         'd2836: data <= 32'h00279793;         'd2837: data <= 32'hff040693;
         'd2838: data <= 32'h00f687b3;         'd2839: data <= 32'hfce7aa23;
         'd2840: data <= 32'hfec42783;         'd2841: data <= 32'h00178793;
         'd2842: data <= 32'hfef42623;         'd2843: data <= 32'hfec42703;
         'd2844: data <= 32'h00700793;         'd2845: data <= 32'hfae7f8e3;
         'd2846: data <= 32'h0480006f;         'd2847: data <= 32'hfa440713;
         'd2848: data <= 32'hfa040793;         'd2849: data <= 32'h00070593;
         'd2850: data <= 32'h00078513;         'd2851: data <= 32'h4b4000ef;
         'd2852: data <= 32'hfea42223;         'd2853: data <= 32'hfe442783;
         'd2854: data <= 32'h00279793;         'd2855: data <= 32'hff040713;
         'd2856: data <= 32'h00f707b3;         'd2857: data <= 32'hfd47a783;
         'd2858: data <= 32'h00178713;         'd2859: data <= 32'hfe442783;
         'd2860: data <= 32'h00279793;         'd2861: data <= 32'hff040693;
         'd2862: data <= 32'h00f687b3;         'd2863: data <= 32'hfce7aa23;
         'd2864: data <= 32'hfa042783;         'd2865: data <= 32'h0007c783;
         'd2866: data <= 32'hfa079ae3;         'd2867: data <= 32'hf9842783;
         'd2868: data <= 32'hfaf42023;         'd2869: data <= 32'h0440006f;
         'd2870: data <= 32'hfa042783;         'd2871: data <= 32'h0007c703;
         'd2872: data <= 32'h02c00793;         'd2873: data <= 32'h02f70263;
         'd2874: data <= 32'hfa042783;         'd2875: data <= 32'h0007c683;
         'd2876: data <= 32'hf9645783;         'd2877: data <= 32'h0ff7f713;
         'd2878: data <= 32'hfa042783;         'd2879: data <= 32'h00e6c733;
         'd2880: data <= 32'h0ff77713;         'd2881: data <= 32'h00e78023;
         'd2882: data <= 32'hfa042703;         'd2883: data <= 32'hf9241783;
         'd2884: data <= 32'h00f707b3;         'd2885: data <= 32'hfaf42023;
         'd2886: data <= 32'hf9842703;         'd2887: data <= 32'hf9c42783;
         'd2888: data <= 32'h00f70733;         'd2889: data <= 32'hfa042783;
         'd2890: data <= 32'hfae7e8e3;         'd2891: data <= 32'hf9842783;
         'd2892: data <= 32'hfaf42023;         'd2893: data <= 32'h0480006f;
         'd2894: data <= 32'hfa440713;         'd2895: data <= 32'hfa040793;
         'd2896: data <= 32'h00070593;         'd2897: data <= 32'h00078513;
         'd2898: data <= 32'h3f8000ef;         'd2899: data <= 32'hfea42423;
         'd2900: data <= 32'hfe842783;         'd2901: data <= 32'h00279793;
         'd2902: data <= 32'hff040713;         'd2903: data <= 32'h00f707b3;
         'd2904: data <= 32'hfd47a783;         'd2905: data <= 32'h00178713;
         'd2906: data <= 32'hfe842783;         'd2907: data <= 32'h00279793;
         'd2908: data <= 32'hff040693;         'd2909: data <= 32'h00f687b3;
         'd2910: data <= 32'hfce7aa23;         'd2911: data <= 32'hfa042783;
         'd2912: data <= 32'h0007c783;         'd2913: data <= 32'hfa079ae3;
         'd2914: data <= 32'hf9842783;         'd2915: data <= 32'hfaf42023;
         'd2916: data <= 32'h0440006f;         'd2917: data <= 32'hfa042783;
         'd2918: data <= 32'h0007c703;         'd2919: data <= 32'h02c00793;
         'd2920: data <= 32'h02f70263;         'd2921: data <= 32'hfa042783;
         'd2922: data <= 32'h0007c683;         'd2923: data <= 32'hf9445783;
         'd2924: data <= 32'h0ff7f713;         'd2925: data <= 32'hfa042783;
         'd2926: data <= 32'h00e6c733;         'd2927: data <= 32'h0ff77713;
         'd2928: data <= 32'h00e78023;         'd2929: data <= 32'hfa042703;
         'd2930: data <= 32'hf9241783;         'd2931: data <= 32'h00f707b3;
         'd2932: data <= 32'hfaf42023;         'd2933: data <= 32'hf9842703;
         'd2934: data <= 32'hf9c42783;         'd2935: data <= 32'h00f70733;
         'd2936: data <= 32'hfa042783;         'd2937: data <= 32'hfae7e8e3;
         'd2938: data <= 32'hfe042623;         'd2939: data <= 32'h0680006f;
         'd2940: data <= 32'hfec42783;         'd2941: data <= 32'h00279793;
         'd2942: data <= 32'hff040713;         'd2943: data <= 32'h00f707b3;
         'd2944: data <= 32'hfd47a783;         'd2945: data <= 32'hf9045703;
         'd2946: data <= 32'h00070593;         'd2947: data <= 32'h00078513;
         'd2948: data <= 32'h0e5000ef;         'd2949: data <= 32'h00050793;
         'd2950: data <= 32'hf8f41823;         'd2951: data <= 32'hfec42783;
         'd2952: data <= 32'h00279793;         'd2953: data <= 32'hff040713;
         'd2954: data <= 32'h00f707b3;         'd2955: data <= 32'hfb47a783;
         'd2956: data <= 32'hf9045703;         'd2957: data <= 32'h00070593;
         'd2958: data <= 32'h00078513;         'd2959: data <= 32'h0b9000ef;
         'd2960: data <= 32'h00050793;         'd2961: data <= 32'hf8f41823;
         'd2962: data <= 32'hfec42783;         'd2963: data <= 32'h00178793;
         'd2964: data <= 32'hfef42623;         'd2965: data <= 32'hfec42703;
         'd2966: data <= 32'h00700793;         'd2967: data <= 32'hf8e7fae3;
         'd2968: data <= 32'hf9045783;         'd2969: data <= 32'h00078513;
         'd2970: data <= 32'h06c12083;         'd2971: data <= 32'h06812403;
         'd2972: data <= 32'h07010113;         'd2973: data <= 32'h00008067;
         'd2974: data <= 32'hfd010113;         'd2975: data <= 32'h02812623;
         'd2976: data <= 32'h03010413;         'd2977: data <= 32'hfca42e23;
         'd2978: data <= 32'h00058793;         'd2979: data <= 32'hfcc42a23;
         'd2980: data <= 32'hfcf41d23;         'd2981: data <= 32'hfe042623;
         'd2982: data <= 32'hfe042423;         'd2983: data <= 32'hfe042023;
         'd2984: data <= 32'hfdc42783;         'd2985: data <= 32'hfff78793;
         'd2986: data <= 32'hfcf42e23;         'd2987: data <= 32'hfe042423;
         'd2988: data <= 32'h1dc0006f;         'd2989: data <= 32'hfe842783;
         'd2990: data <= 32'h06078e63;         'd2991: data <= 32'hfe042223;
         'd2992: data <= 32'h0380006f;         'd2993: data <= 32'hfe042703;
         'd2994: data <= 32'hfe442783;         'd2995: data <= 32'h00f70733;
         'd2996: data <= 32'hfec42683;         'd2997: data <= 32'hfe442783;
         'd2998: data <= 32'h00f687b3;         'd2999: data <= 32'hfd442683;
         'd3000: data <= 32'h00f687b3;         'd3001: data <= 32'h00074703;
         'd3002: data <= 32'h00e78023;         'd3003: data <= 32'hfe442783;
         'd3004: data <= 32'h00178793;         'd3005: data <= 32'hfef42223;
         'd3006: data <= 32'hfe442703;         'd3007: data <= 32'hfe842783;
         'd3008: data <= 32'hfcf762e3;         'd3009: data <= 32'hfec42703;
         'd3010: data <= 32'hfe442783;         'd3011: data <= 32'h00f707b3;
         'd3012: data <= 32'hfd442703;         'd3013: data <= 32'h00f707b3;
         'd3014: data <= 32'h02c00713;         'd3015: data <= 32'h00e78023;
         'd3016: data <= 32'hfe842703;         'd3017: data <= 32'hfec42783;
         'd3018: data <= 32'h00f707b3;         'd3019: data <= 32'h00178793;
         'd3020: data <= 32'hfef42623;         'd3021: data <= 32'hfda41783;
         'd3022: data <= 32'h01079793;         'd3023: data <= 32'h0107d793;
         'd3024: data <= 32'h00178793;         'd3025: data <= 32'h01079793;
         'd3026: data <= 32'h0107d793;         'd3027: data <= 32'hfcf41d23;
         'd3028: data <= 32'hfda45783;         'd3029: data <= 32'h0077f793;
         'd3030: data <= 32'h00700713;         'd3031: data <= 32'h0ee78863;
         'd3032: data <= 32'h00700713;         'd3033: data <= 32'h12f74263;
         'd3034: data <= 32'h00600713;         'd3035: data <= 32'h10f74e63;
         'd3036: data <= 32'h00500713;         'd3037: data <= 32'h08e7de63;
         'd3038: data <= 32'h00200713;         'd3039: data <= 32'h00f74663;
         'd3040: data <= 32'h0007dc63;         'd3041: data <= 32'h1040006f;
         'd3042: data <= 32'hffd78713;         'd3043: data <= 32'h00100793;
         'd3044: data <= 32'h0ee7ec63;         'd3045: data <= 32'h0400006f;
         'd3046: data <= 32'hfda41783;         'd3047: data <= 32'h4037d793;
         'd3048: data <= 32'h01079793;         'd3049: data <= 32'h4107d793;
         'd3050: data <= 32'h01079793;         'd3051: data <= 32'h0107d793;
         'd3052: data <= 32'h0037f793;         'd3053: data <= 32'h83018713;
         'd3054: data <= 32'h00279793;         'd3055: data <= 32'h00f707b3;
         'd3056: data <= 32'h0007a783;         'd3057: data <= 32'hfef42023;
         'd3058: data <= 32'h00400793;         'd3059: data <= 32'hfef42423;
         'd3060: data <= 32'h0bc0006f;         'd3061: data <= 32'hfda41783;
         'd3062: data <= 32'h4037d793;         'd3063: data <= 32'h01079793;
         'd3064: data <= 32'h4107d793;         'd3065: data <= 32'h01079793;
         'd3066: data <= 32'h0107d793;         'd3067: data <= 32'h0037f793;
         'd3068: data <= 32'h84018713;         'd3069: data <= 32'h00279793;
         'd3070: data <= 32'h00f707b3;         'd3071: data <= 32'h0007a783;
         'd3072: data <= 32'hfef42023;         'd3073: data <= 32'h00800793;
         'd3074: data <= 32'hfef42423;         'd3075: data <= 32'h0800006f;
         'd3076: data <= 32'hfda41783;         'd3077: data <= 32'h4037d793;
         'd3078: data <= 32'h01079793;         'd3079: data <= 32'h4107d793;
         'd3080: data <= 32'h01079793;         'd3081: data <= 32'h0107d793;
         'd3082: data <= 32'h0037f793;         'd3083: data <= 32'h85018713;
         'd3084: data <= 32'h00279793;         'd3085: data <= 32'h00f707b3;
         'd3086: data <= 32'h0007a783;         'd3087: data <= 32'hfef42023;
         'd3088: data <= 32'h00800793;         'd3089: data <= 32'hfef42423;
         'd3090: data <= 32'h0440006f;         'd3091: data <= 32'hfda41783;
         'd3092: data <= 32'h4037d793;         'd3093: data <= 32'h01079793;
         'd3094: data <= 32'h4107d793;         'd3095: data <= 32'h01079793;
         'd3096: data <= 32'h0107d793;         'd3097: data <= 32'h0037f793;
         'd3098: data <= 32'h86018713;         'd3099: data <= 32'h00279793;
         'd3100: data <= 32'h00f707b3;         'd3101: data <= 32'h0007a783;
         'd3102: data <= 32'hfef42023;         'd3103: data <= 32'h00800793;
         'd3104: data <= 32'hfef42423;         'd3105: data <= 32'h0080006f;
         'd3106: data <= 32'h00000013;         'd3107: data <= 32'hfec42703;
         'd3108: data <= 32'hfe842783;         'd3109: data <= 32'h00f707b3;
         'd3110: data <= 32'h00178793;         'd3111: data <= 32'hfdc42703;
         'd3112: data <= 32'he0e7eae3;         'd3113: data <= 32'hfdc42783;
         'd3114: data <= 32'h00178793;         'd3115: data <= 32'hfcf42e23;
         'd3116: data <= 32'h0200006f;         'd3117: data <= 32'hfd442703;
         'd3118: data <= 32'hfec42783;         'd3119: data <= 32'h00f707b3;
         'd3120: data <= 32'h00078023;         'd3121: data <= 32'hfec42783;
         'd3122: data <= 32'h00178793;         'd3123: data <= 32'hfef42623;
         'd3124: data <= 32'hfec42703;         'd3125: data <= 32'hfdc42783;
         'd3126: data <= 32'hfcf76ee3;         'd3127: data <= 32'h00000013;
         'd3128: data <= 32'h00000013;         'd3129: data <= 32'h02c12403;
         'd3130: data <= 32'h03010113;         'd3131: data <= 32'h00008067;
         'd3132: data <= 32'hfd010113;         'd3133: data <= 32'h02812623;
         'd3134: data <= 32'h03010413;         'd3135: data <= 32'h00050793;
         'd3136: data <= 32'hfcf40fa3;         'd3137: data <= 32'hfdf44783;
         'd3138: data <= 32'h0307b793;         'd3139: data <= 32'h0017c793;
         'd3140: data <= 32'h0ff7f713;         'd3141: data <= 32'hfdf44783;
         'd3142: data <= 32'h03a7b793;         'd3143: data <= 32'h0ff7f793;
         'd3144: data <= 32'h00f777b3;         'd3145: data <= 32'h0ff7f793;
         'd3146: data <= 32'hfef407a3;         'd3147: data <= 32'hfef44783;
         'd3148: data <= 32'h00078513;         'd3149: data <= 32'h02c12403;
         'd3150: data <= 32'h03010113;         'd3151: data <= 32'h00008067;
         'd3152: data <= 32'hfd010113;         'd3153: data <= 32'h02112623;
         'd3154: data <= 32'h02812423;         'd3155: data <= 32'h03010413;
         'd3156: data <= 32'hfca42e23;         'd3157: data <= 32'hfcb42c23;
         'd3158: data <= 32'hfdc42783;         'd3159: data <= 32'h0007a783;
         'd3160: data <= 32'hfef42623;         'd3161: data <= 32'hfe042423;
         'd3162: data <= 32'h3380006f;         'd3163: data <= 32'hfec42783;
         'd3164: data <= 32'h0007c783;         'd3165: data <= 32'hfef403a3;
         'd3166: data <= 32'hfe744703;         'd3167: data <= 32'h02c00793;
         'd3168: data <= 32'h00f71a63;         'd3169: data <= 32'hfec42783;
         'd3170: data <= 32'h00178793;         'd3171: data <= 32'hfef42623;
         'd3172: data <= 32'h3280006f;         'd3173: data <= 32'hfe842703;
         'd3174: data <= 32'h00700793;         'd3175: data <= 32'h2ce7ee63;
         'd3176: data <= 32'hfe842783;         'd3177: data <= 32'h00279713;
         'd3178: data <= 32'h800057b7;         'd3179: data <= 32'h5d078793;
         'd3180: data <= 32'h00f707b3;         'd3181: data <= 32'h0007a783;
         'd3182: data <= 32'h00078067;         'd3183: data <= 32'hfe744783;
         'd3184: data <= 32'h00078513;         'd3185: data <= 32'hf2dff0ef;
         'd3186: data <= 32'h00050793;         'd3187: data <= 32'h00078863;
         'd3188: data <= 32'h00400793;         'd3189: data <= 32'hfef42423;
         'd3190: data <= 32'h05c0006f;         'd3191: data <= 32'hfe744703;
         'd3192: data <= 32'h02b00793;         'd3193: data <= 32'h00f70863;
         'd3194: data <= 32'hfe744703;         'd3195: data <= 32'h02d00793;
         'd3196: data <= 32'h00f71863;         'd3197: data <= 32'h00200793;
         'd3198: data <= 32'hfef42423;         'd3199: data <= 32'h0380006f;
         'd3200: data <= 32'hfe744703;         'd3201: data <= 32'h02e00793;
         'd3202: data <= 32'h00f71863;         'd3203: data <= 32'h00500793;
         'd3204: data <= 32'hfef42423;         'd3205: data <= 32'h0200006f;
         'd3206: data <= 32'h00100793;         'd3207: data <= 32'hfef42423;
         'd3208: data <= 32'hfd842783;         'd3209: data <= 32'h00478793;
         'd3210: data <= 32'h0007a703;         'd3211: data <= 32'h00170713;
         'd3212: data <= 32'h00e7a023;         'd3213: data <= 32'hfd842783;
         'd3214: data <= 32'h0007a783;         'd3215: data <= 32'h00178713;
         'd3216: data <= 32'hfd842783;         'd3217: data <= 32'h00e7a023;
         'd3218: data <= 32'h24c0006f;         'd3219: data <= 32'hfe744783;
         'd3220: data <= 32'h00078513;         'd3221: data <= 32'he9dff0ef;
         'd3222: data <= 32'h00050793;         'd3223: data <= 32'h02078263;
         'd3224: data <= 32'h00400793;         'd3225: data <= 32'hfef42423;
         'd3226: data <= 32'hfd842783;         'd3227: data <= 32'h00878793;
         'd3228: data <= 32'h0007a703;         'd3229: data <= 32'h00170713;
         'd3230: data <= 32'h00e7a023;         'd3231: data <= 32'h2180006f;
         'd3232: data <= 32'hfe744703;         'd3233: data <= 32'h02e00793;
         'd3234: data <= 32'h02f71263;         'd3235: data <= 32'h00500793;
         'd3236: data <= 32'hfef42423;         'd3237: data <= 32'hfd842783;
         'd3238: data <= 32'h00878793;         'd3239: data <= 32'h0007a703;
         'd3240: data <= 32'h00170713;         'd3241: data <= 32'h00e7a023;
         'd3242: data <= 32'h1ec0006f;         'd3243: data <= 32'h00100793;
         'd3244: data <= 32'hfef42423;         'd3245: data <= 32'hfd842783;
         'd3246: data <= 32'h00878793;         'd3247: data <= 32'h0007a703;
         'd3248: data <= 32'h00170713;         'd3249: data <= 32'h00e7a023;
         'd3250: data <= 32'h1cc0006f;         'd3251: data <= 32'hfe744703;
         'd3252: data <= 32'h02e00793;         'd3253: data <= 32'h02f71263;
         'd3254: data <= 32'h00500793;         'd3255: data <= 32'hfef42423;
         'd3256: data <= 32'hfd842783;         'd3257: data <= 32'h01078793;
         'd3258: data <= 32'h0007a703;         'd3259: data <= 32'h00170713;
         'd3260: data <= 32'h00e7a023;         'd3261: data <= 32'h18c0006f;
         'd3262: data <= 32'hfe744783;         'd3263: data <= 32'h00078513;
         'd3264: data <= 32'hdf1ff0ef;         'd3265: data <= 32'h00050793;
         'd3266: data <= 32'h16079c63;         'd3267: data <= 32'h00100793;
         'd3268: data <= 32'hfef42423;         'd3269: data <= 32'hfd842783;
         'd3270: data <= 32'h01078793;         'd3271: data <= 32'h0007a703;
         'd3272: data <= 32'h00170713;         'd3273: data <= 32'h00e7a023;
         'd3274: data <= 32'h1580006f;         'd3275: data <= 32'hfe744703;
         'd3276: data <= 32'h04500793;         'd3277: data <= 32'h00f70863;
         'd3278: data <= 32'hfe744703;         'd3279: data <= 32'h06500793;
         'd3280: data <= 32'h02f71263;         'd3281: data <= 32'h00300793;
         'd3282: data <= 32'hfef42423;         'd3283: data <= 32'hfd842783;
         'd3284: data <= 32'h01478793;         'd3285: data <= 32'h0007a703;
         'd3286: data <= 32'h00170713;         'd3287: data <= 32'h00e7a023;
         'd3288: data <= 32'h1280006f;         'd3289: data <= 32'hfe744783;
         'd3290: data <= 32'h00078513;         'd3291: data <= 32'hd85ff0ef;
         'd3292: data <= 32'h00050793;         'd3293: data <= 32'h10079a63;
         'd3294: data <= 32'h00100793;         'd3295: data <= 32'hfef42423;
         'd3296: data <= 32'hfd842783;         'd3297: data <= 32'h01478793;
         'd3298: data <= 32'h0007a703;         'd3299: data <= 32'h00170713;
         'd3300: data <= 32'h00e7a023;         'd3301: data <= 32'h0f40006f;
         'd3302: data <= 32'hfe744703;         'd3303: data <= 32'h02b00793;
         'd3304: data <= 32'h00f70863;         'd3305: data <= 32'hfe744703;
         'd3306: data <= 32'h02d00793;         'd3307: data <= 32'h02f71263;
         'd3308: data <= 32'h00600793;         'd3309: data <= 32'hfef42423;
         'd3310: data <= 32'hfd842783;         'd3311: data <= 32'h00c78793;
         'd3312: data <= 32'h0007a703;         'd3313: data <= 32'h00170713;
         'd3314: data <= 32'h00e7a023;         'd3315: data <= 32'h0c80006f;
         'd3316: data <= 32'h00100793;         'd3317: data <= 32'hfef42423;
         'd3318: data <= 32'hfd842783;         'd3319: data <= 32'h00c78793;
         'd3320: data <= 32'h0007a703;         'd3321: data <= 32'h00170713;
         'd3322: data <= 32'h00e7a023;         'd3323: data <= 32'h0a80006f;
         'd3324: data <= 32'hfe744783;         'd3325: data <= 32'h00078513;
         'd3326: data <= 32'hcf9ff0ef;         'd3327: data <= 32'h00050793;
         'd3328: data <= 32'h02078263;         'd3329: data <= 32'h00700793;
         'd3330: data <= 32'hfef42423;         'd3331: data <= 32'hfd842783;
         'd3332: data <= 32'h01878793;         'd3333: data <= 32'h0007a703;
         'd3334: data <= 32'h00170713;         'd3335: data <= 32'h00e7a023;
         'd3336: data <= 32'h0740006f;         'd3337: data <= 32'h00100793;
         'd3338: data <= 32'hfef42423;         'd3339: data <= 32'hfd842783;
         'd3340: data <= 32'h01878793;         'd3341: data <= 32'h0007a703;
         'd3342: data <= 32'h00170713;         'd3343: data <= 32'h00e7a023;
         'd3344: data <= 32'h0540006f;         'd3345: data <= 32'hfe744783;
         'd3346: data <= 32'h00078513;         'd3347: data <= 32'hca5ff0ef;
         'd3348: data <= 32'h00050793;         'd3349: data <= 32'h02079e63;
         'd3350: data <= 32'h00100793;         'd3351: data <= 32'hfef42423;
         'd3352: data <= 32'hfd842783;         'd3353: data <= 32'h00478793;
         'd3354: data <= 32'h0007a703;         'd3355: data <= 32'h00170713;
         'd3356: data <= 32'h00e7a023;         'd3357: data <= 32'h01c0006f;
         'd3358: data <= 32'h00000013;         'd3359: data <= 32'h0180006f;
         'd3360: data <= 32'h00000013;         'd3361: data <= 32'h0100006f;
         'd3362: data <= 32'h00000013;         'd3363: data <= 32'h0080006f;
         'd3364: data <= 32'h00000013;         'd3365: data <= 32'hfec42783;
         'd3366: data <= 32'h00178793;         'd3367: data <= 32'hfef42623;
         'd3368: data <= 32'hfec42783;         'd3369: data <= 32'h0007c783;
         'd3370: data <= 32'h00078863;         'd3371: data <= 32'hfe842703;
         'd3372: data <= 32'h00100793;         'd3373: data <= 32'hcaf71ce3;
         'd3374: data <= 32'hfdc42783;         'd3375: data <= 32'hfec42703;
         'd3376: data <= 32'h00e7a023;         'd3377: data <= 32'hfe842783;
         'd3378: data <= 32'h00078513;         'd3379: data <= 32'h02c12083;
         'd3380: data <= 32'h02812403;         'd3381: data <= 32'h03010113;
         'd3382: data <= 32'h00008067;         'd3383: data <= 32'hfd010113;
         'd3384: data <= 32'h02812623;         'd3385: data <= 32'h03010413;
         'd3386: data <= 32'hfca42e23;         'd3387: data <= 32'hfdc42703;
         'd3388: data <= 32'h00500793;         'd3389: data <= 32'h04e7ee63;
         'd3390: data <= 32'hfdc42783;         'd3391: data <= 32'h00279713;
         'd3392: data <= 32'h800057b7;         'd3393: data <= 32'h5f078793;
         'd3394: data <= 32'h00f707b3;         'd3395: data <= 32'h0007a783;
         'd3396: data <= 32'h00078067;         'd3397: data <= 32'h8801a783;
         'd3398: data <= 32'hfef42623;         'd3399: data <= 32'h03c0006f;
         'd3400: data <= 32'h8841a783;         'd3401: data <= 32'hfef42623;
         'd3402: data <= 32'h0300006f;         'd3403: data <= 32'h8701a783;
         'd3404: data <= 32'hfef42623;         'd3405: data <= 32'h0240006f;
         'd3406: data <= 32'h8881a783;         'd3407: data <= 32'hfef42623;
         'd3408: data <= 32'h0180006f;         'd3409: data <= 32'h88c1a783;
         'd3410: data <= 32'hfef42623;         'd3411: data <= 32'h00c0006f;
         'd3412: data <= 32'hfe042623;         'd3413: data <= 32'h00000013;
         'd3414: data <= 32'hfec42783;         'd3415: data <= 32'h00078513;
         'd3416: data <= 32'h02c12403;         'd3417: data <= 32'h03010113;
         'd3418: data <= 32'h00008067;         'd3419: data <= 32'hfd010113;
         'd3420: data <= 32'h02812623;         'd3421: data <= 32'h03010413;
         'd3422: data <= 32'h00050793;         'd3423: data <= 32'h00058713;
         'd3424: data <= 32'hfcf40fa3;         'd3425: data <= 32'h00070793;
         'd3426: data <= 32'hfcf41e23;         'd3427: data <= 32'hfe0407a3;
         'd3428: data <= 32'hfe0406a3;         'd3429: data <= 32'hfe040723;
         'd3430: data <= 32'hfe0407a3;         'd3431: data <= 32'h0b00006f;
         'd3432: data <= 32'hfdc45783;         'd3433: data <= 32'h01879713;
         'd3434: data <= 32'h41875713;         'd3435: data <= 32'hfdf40783;
         'd3436: data <= 32'h00f747b3;         'd3437: data <= 32'h01879793;
         'd3438: data <= 32'h4187d793;         'd3439: data <= 32'h0ff7f793;
         'd3440: data <= 32'h0017f793;         'd3441: data <= 32'hfef406a3;
         'd3442: data <= 32'hfdf44783;         'd3443: data <= 32'h0017d793;
         'd3444: data <= 32'hfcf40fa3;         'd3445: data <= 32'hfed44703;
         'd3446: data <= 32'h00100793;         'd3447: data <= 32'h02f71263;
         'd3448: data <= 32'hfdc45703;         'd3449: data <= 32'h000047b7;
         'd3450: data <= 32'h00278793;         'd3451: data <= 32'h00f747b3;
         'd3452: data <= 32'hfcf41e23;         'd3453: data <= 32'h00100793;
         'd3454: data <= 32'hfef40723;         'd3455: data <= 32'h0080006f;
         'd3456: data <= 32'hfe040723;         'd3457: data <= 32'hfdc45783;
         'd3458: data <= 32'h0017d793;         'd3459: data <= 32'hfcf41e23;
         'd3460: data <= 32'hfee44783;         'd3461: data <= 32'h00078c63;
         'd3462: data <= 32'hfdc45703;         'd3463: data <= 32'hffff87b7;
         'd3464: data <= 32'h00f767b3;         'd3465: data <= 32'hfcf41e23;
         'd3466: data <= 32'h0180006f;         'd3467: data <= 32'hfdc45703;
         'd3468: data <= 32'h000087b7;         'd3469: data <= 32'hfff78793;
         'd3470: data <= 32'h00f777b3;         'd3471: data <= 32'hfcf41e23;
         'd3472: data <= 32'hfef44783;         'd3473: data <= 32'h00178793;
         'd3474: data <= 32'hfef407a3;         'd3475: data <= 32'hfef44703;
         'd3476: data <= 32'h00700793;         'd3477: data <= 32'hf4e7f6e3;
         'd3478: data <= 32'hfdc45783;         'd3479: data <= 32'h00078513;
         'd3480: data <= 32'h02c12403;         'd3481: data <= 32'h03010113;
         'd3482: data <= 32'h00008067;         'd3483: data <= 32'hfe010113;
         'd3484: data <= 32'h00112e23;         'd3485: data <= 32'h00812c23;
         'd3486: data <= 32'h02010413;         'd3487: data <= 32'h00050793;
         'd3488: data <= 32'h00058713;         'd3489: data <= 32'hfef41723;
         'd3490: data <= 32'h00070793;         'd3491: data <= 32'hfef41623;
         'd3492: data <= 32'hfee45783;         'd3493: data <= 32'h0ff7f793;
         'd3494: data <= 32'hfec45703;         'd3495: data <= 32'h00070593;
         'd3496: data <= 32'h00078513;         'd3497: data <= 32'hec9ff0ef;
         'd3498: data <= 32'h00050793;         'd3499: data <= 32'hfef41623;
         'd3500: data <= 32'hfee45783;         'd3501: data <= 32'h0087d793;
         'd3502: data <= 32'h01079793;         'd3503: data <= 32'h0107d793;
         'd3504: data <= 32'h0ff7f793;         'd3505: data <= 32'hfec45703;
         'd3506: data <= 32'h00070593;         'd3507: data <= 32'h00078513;
         'd3508: data <= 32'he9dff0ef;         'd3509: data <= 32'h00050793;
         'd3510: data <= 32'hfef41623;         'd3511: data <= 32'hfec45783;
         'd3512: data <= 32'h00078513;         'd3513: data <= 32'h01c12083;
         'd3514: data <= 32'h01812403;         'd3515: data <= 32'h02010113;
         'd3516: data <= 32'h00008067;         'd3517: data <= 32'hfe010113;
         'd3518: data <= 32'h00112e23;         'd3519: data <= 32'h00812c23;
         'd3520: data <= 32'h02010413;         'd3521: data <= 32'hfea42623;
         'd3522: data <= 32'h00058793;         'd3523: data <= 32'hfef41523;
         'd3524: data <= 32'hfec42783;         'd3525: data <= 32'h01079793;
         'd3526: data <= 32'h4107d793;         'd3527: data <= 32'hfea45703;
         'd3528: data <= 32'h00070593;         'd3529: data <= 32'h00078513;
         'd3530: data <= 32'h04c000ef;         'd3531: data <= 32'h00050793;
         'd3532: data <= 32'hfef41523;         'd3533: data <= 32'hfec42783;
         'd3534: data <= 32'h0107d793;         'd3535: data <= 32'h01079793;
         'd3536: data <= 32'h4107d793;         'd3537: data <= 32'hfea45703;
         'd3538: data <= 32'h00070593;         'd3539: data <= 32'h00078513;
         'd3540: data <= 32'h024000ef;         'd3541: data <= 32'h00050793;
         'd3542: data <= 32'hfef41523;         'd3543: data <= 32'hfea45783;
         'd3544: data <= 32'h00078513;         'd3545: data <= 32'h01c12083;
         'd3546: data <= 32'h01812403;         'd3547: data <= 32'h02010113;
         'd3548: data <= 32'h00008067;         'd3549: data <= 32'hfe010113;
         'd3550: data <= 32'h00112e23;         'd3551: data <= 32'h00812c23;
         'd3552: data <= 32'h02010413;         'd3553: data <= 32'h00050793;
         'd3554: data <= 32'h00058713;         'd3555: data <= 32'hfef41723;
         'd3556: data <= 32'h00070793;         'd3557: data <= 32'hfef41623;
         'd3558: data <= 32'hfee45783;         'd3559: data <= 32'hfec45703;
         'd3560: data <= 32'h00070593;         'd3561: data <= 32'h00078513;
         'd3562: data <= 32'hec5ff0ef;         'd3563: data <= 32'h00050793;
         'd3564: data <= 32'h00078513;         'd3565: data <= 32'h01c12083;
         'd3566: data <= 32'h01812403;         'd3567: data <= 32'h02010113;
         'd3568: data <= 32'h00008067;         'd3569: data <= 32'hfe010113;
         'd3570: data <= 32'h00112e23;         'd3571: data <= 32'h00812c23;
         'd3572: data <= 32'h02010413;         'd3573: data <= 32'hfe0407a3;
         'd3574: data <= 32'hfef44783;         'd3575: data <= 32'h00078863;
         'd3576: data <= 32'h800057b7;         'd3577: data <= 32'h60878513;
         'd3578: data <= 32'h2b8010ef;         'd3579: data <= 32'hfef44783;
         'd3580: data <= 32'h00078513;         'd3581: data <= 32'h01c12083;
         'd3582: data <= 32'h01812403;         'd3583: data <= 32'h02010113;
         'd3584: data <= 32'h00008067;         'd3585: data <= 32'hfe010113;
         'd3586: data <= 32'h00812e23;         'd3587: data <= 32'h02010413;
         'd3588: data <= 32'h00050793;         'd3589: data <= 32'hfeb42423;
         'd3590: data <= 32'hfec42223;         'd3591: data <= 32'hfed42023;
         'd3592: data <= 32'hfef407a3;         'd3593: data <= 32'hfe442703;
         'd3594: data <= 32'hfe042783;         'd3595: data <= 32'h00f77c63;
         'd3596: data <= 32'hfe842703;         'd3597: data <= 32'hfe442783;
         'd3598: data <= 32'h00f707b3;         'd3599: data <= 32'hfef44703;
         'd3600: data <= 32'h00e78023;         'd3601: data <= 32'h00000013;
         'd3602: data <= 32'h01c12403;         'd3603: data <= 32'h02010113;
         'd3604: data <= 32'h00008067;         'd3605: data <= 32'hfe010113;
         'd3606: data <= 32'h00812e23;         'd3607: data <= 32'h02010413;
         'd3608: data <= 32'h00050793;         'd3609: data <= 32'hfeb42423;
         'd3610: data <= 32'hfec42223;         'd3611: data <= 32'hfed42023;
         'd3612: data <= 32'hfef407a3;         'd3613: data <= 32'h00000013;
         'd3614: data <= 32'h01c12403;         'd3615: data <= 32'h02010113;
         'd3616: data <= 32'h00008067;         'd3617: data <= 32'hfe010113;
         'd3618: data <= 32'h00112e23;         'd3619: data <= 32'h00812c23;
         'd3620: data <= 32'h02010413;         'd3621: data <= 32'h00050793;
         'd3622: data <= 32'hfeb42423;         'd3623: data <= 32'hfec42223;
         'd3624: data <= 32'hfed42023;         'd3625: data <= 32'hfef407a3;
         'd3626: data <= 32'hfef44783;         'd3627: data <= 32'h00078863;
         'd3628: data <= 32'hfef44783;         'd3629: data <= 32'h00078513;
         'd3630: data <= 32'h49c010ef;         'd3631: data <= 32'h00000013;
         'd3632: data <= 32'h01c12083;         'd3633: data <= 32'h01812403;
         'd3634: data <= 32'h02010113;         'd3635: data <= 32'h00008067;
         'd3636: data <= 32'hfe010113;         'd3637: data <= 32'h00112e23;
         'd3638: data <= 32'h00812c23;         'd3639: data <= 32'h02010413;
         'd3640: data <= 32'h00050793;         'd3641: data <= 32'hfeb42423;
         'd3642: data <= 32'hfec42223;         'd3643: data <= 32'hfed42023;
         'd3644: data <= 32'hfef407a3;         'd3645: data <= 32'hfef44783;
         'd3646: data <= 32'h02078263;         'd3647: data <= 32'hfe842783;
         'd3648: data <= 32'h0007a683;         'd3649: data <= 32'hfe842783;
         'd3650: data <= 32'h0047a703;         'd3651: data <= 32'hfef44783;
         'd3652: data <= 32'h00070593;         'd3653: data <= 32'h00078513;
         'd3654: data <= 32'h000680e7;         'd3655: data <= 32'h00000013;
         'd3656: data <= 32'h01c12083;         'd3657: data <= 32'h01812403;
         'd3658: data <= 32'h02010113;         'd3659: data <= 32'h00008067;
         'd3660: data <= 32'hfd010113;         'd3661: data <= 32'h02812623;
         'd3662: data <= 32'h03010413;         'd3663: data <= 32'hfca42e23;
         'd3664: data <= 32'hfcb42c23;         'd3665: data <= 32'hfdc42783;
         'd3666: data <= 32'hfef42623;         'd3667: data <= 32'h0100006f;
         'd3668: data <= 32'hfec42783;         'd3669: data <= 32'h00178793;
         'd3670: data <= 32'hfef42623;         'd3671: data <= 32'hfec42783;
         'd3672: data <= 32'h0007c783;         'd3673: data <= 32'h00078a63;
         'd3674: data <= 32'hfd842783;         'd3675: data <= 32'hfff78713;
         'd3676: data <= 32'hfce42c23;         'd3677: data <= 32'hfc079ee3;
         'd3678: data <= 32'hfec42703;         'd3679: data <= 32'hfdc42783;
         'd3680: data <= 32'h40f707b3;         'd3681: data <= 32'h00078513;
         'd3682: data <= 32'h02c12403;         'd3683: data <= 32'h03010113;
         'd3684: data <= 32'h00008067;         'd3685: data <= 32'hfe010113;
         'd3686: data <= 32'h00812e23;         'd3687: data <= 32'h02010413;
         'd3688: data <= 32'h00050793;         'd3689: data <= 32'hfef407a3;
         'd3690: data <= 32'hfef44703;         'd3691: data <= 32'h02f00793;
         'd3692: data <= 32'h00e7fc63;         'd3693: data <= 32'hfef44703;
         'd3694: data <= 32'h03900793;         'd3695: data <= 32'h00e7e663;
         'd3696: data <= 32'h00100793;         'd3697: data <= 32'h0080006f;
         'd3698: data <= 32'h00000793;         'd3699: data <= 32'h0017f793;
         'd3700: data <= 32'h0ff7f793;         'd3701: data <= 32'h00078513;
         'd3702: data <= 32'h01c12403;         'd3703: data <= 32'h02010113;
         'd3704: data <= 32'h00008067;         'd3705: data <= 32'hfd010113;
         'd3706: data <= 32'h02112623;         'd3707: data <= 32'h02812423;
         'd3708: data <= 32'h03010413;         'd3709: data <= 32'hfca42e23;
         'd3710: data <= 32'hfe042623;         'd3711: data <= 32'h0400006f;
         'd3712: data <= 32'hfec42703;         'd3713: data <= 32'h00070793;
         'd3714: data <= 32'h00279793;         'd3715: data <= 32'h00e787b3;
         'd3716: data <= 32'h00179793;         'd3717: data <= 32'h00078613;
         'd3718: data <= 32'hfdc42783;         'd3719: data <= 32'h0007a783;
         'd3720: data <= 32'h00178693;         'd3721: data <= 32'hfdc42703;
         'd3722: data <= 32'h00d72023;         'd3723: data <= 32'h0007c783;
         'd3724: data <= 32'h00f607b3;         'd3725: data <= 32'hfd078793;
         'd3726: data <= 32'hfef42623;         'd3727: data <= 32'hfdc42783;
         'd3728: data <= 32'h0007a783;         'd3729: data <= 32'h0007c783;
         'd3730: data <= 32'h00078513;         'd3731: data <= 32'hf49ff0ef;
         'd3732: data <= 32'h00050793;         'd3733: data <= 32'hfa0796e3;
         'd3734: data <= 32'hfec42783;         'd3735: data <= 32'h00078513;
         'd3736: data <= 32'h02c12083;         'd3737: data <= 32'h02812403;
         'd3738: data <= 32'h03010113;         'd3739: data <= 32'h00008067;
         'd3740: data <= 32'hfc010113;         'd3741: data <= 32'h02112e23;
         'd3742: data <= 32'h02812c23;         'd3743: data <= 32'h04010413;
         'd3744: data <= 32'hfca42e23;         'd3745: data <= 32'hfcb42c23;
         'd3746: data <= 32'hfcc42a23;         'd3747: data <= 32'hfcd42823;
         'd3748: data <= 32'hfce42623;         'd3749: data <= 32'hfcf42423;
         'd3750: data <= 32'hfd042223;         'd3751: data <= 32'hfd142023;
         'd3752: data <= 32'hfd442783;         'd3753: data <= 32'hfef42423;
         'd3754: data <= 32'hfc042783;         'd3755: data <= 32'h0027f793;
         'd3756: data <= 32'h08079c63;         'd3757: data <= 32'hfc042783;
         'd3758: data <= 32'h0017f793;         'd3759: data <= 32'h08079663;
         'd3760: data <= 32'hfc842783;         'd3761: data <= 32'hfef42623;
         'd3762: data <= 32'h0340006f;         'd3763: data <= 32'hfd442783;
         'd3764: data <= 32'h00178713;         'd3765: data <= 32'hfce42a23;
         'd3766: data <= 32'hfdc42703;         'd3767: data <= 32'hfd042683;
         'd3768: data <= 32'h00078613;         'd3769: data <= 32'hfd842583;
         'd3770: data <= 32'h02000513;         'd3771: data <= 32'h000700e7;
         'd3772: data <= 32'hfec42783;         'd3773: data <= 32'h00178793;
         'd3774: data <= 32'hfef42623;         'd3775: data <= 32'hfec42703;
         'd3776: data <= 32'hfc442783;         'd3777: data <= 32'hfcf764e3;
         'd3778: data <= 32'h0400006f;         'd3779: data <= 32'hfc842783;
         'd3780: data <= 32'hfff78793;         'd3781: data <= 32'hfcf42423;
         'd3782: data <= 32'hfcc42703;         'd3783: data <= 32'hfc842783;
         'd3784: data <= 32'h00f707b3;         'd3785: data <= 32'h0007c503;
         'd3786: data <= 32'hfd442783;         'd3787: data <= 32'h00178713;
         'd3788: data <= 32'hfce42a23;         'd3789: data <= 32'hfdc42703;
         'd3790: data <= 32'hfd042683;         'd3791: data <= 32'h00078613;
         'd3792: data <= 32'hfd842583;         'd3793: data <= 32'h000700e7;
         'd3794: data <= 32'hfc842783;         'd3795: data <= 32'hfc0790e3;
         'd3796: data <= 32'hfc042783;         'd3797: data <= 32'h0027f793;
         'd3798: data <= 32'h04078063;         'd3799: data <= 32'h0280006f;
         'd3800: data <= 32'hfd442783;         'd3801: data <= 32'h00178713;
         'd3802: data <= 32'hfce42a23;         'd3803: data <= 32'hfdc42703;
         'd3804: data <= 32'hfd042683;         'd3805: data <= 32'h00078613;
         'd3806: data <= 32'hfd842583;         'd3807: data <= 32'h02000513;
         'd3808: data <= 32'h000700e7;         'd3809: data <= 32'hfd442703;
         'd3810: data <= 32'hfe842783;         'd3811: data <= 32'h40f707b3;
         'd3812: data <= 32'hfc442703;         'd3813: data <= 32'hfce7e6e3;
         'd3814: data <= 32'hfd442783;         'd3815: data <= 32'h00078513;
         'd3816: data <= 32'h03c12083;         'd3817: data <= 32'h03812403;
         'd3818: data <= 32'h04010113;         'd3819: data <= 32'h00008067;
         'd3820: data <= 32'hfd010113;         'd3821: data <= 32'h02112623;
         'd3822: data <= 32'h02812423;         'd3823: data <= 32'h03010413;
         'd3824: data <= 32'hfea42623;         'd3825: data <= 32'hfeb42423;
         'd3826: data <= 32'hfec42223;         'd3827: data <= 32'hfed42023;
         'd3828: data <= 32'hfce42e23;         'd3829: data <= 32'hfcf42c23;
         'd3830: data <= 32'h00080793;         'd3831: data <= 32'hfd142823;
         'd3832: data <= 32'hfcf40ba3;         'd3833: data <= 32'h00842783;
         'd3834: data <= 32'h0027f793;         'd3835: data <= 32'h0a079a63;
         'd3836: data <= 32'h00442783;         'd3837: data <= 32'h04078863;
         'd3838: data <= 32'h00842783;         'd3839: data <= 32'h0017f793;
         'd3840: data <= 32'h04078263;         'd3841: data <= 32'hfd744783;
         'd3842: data <= 32'h00079863;         'd3843: data <= 32'h00842783;
         'd3844: data <= 32'h00c7f793;         'd3845: data <= 32'h02078863;
         'd3846: data <= 32'h00442783;         'd3847: data <= 32'hfff78793;
         'd3848: data <= 32'h00f42223;         'd3849: data <= 32'h0200006f;
         'd3850: data <= 32'hfd842783;         'd3851: data <= 32'h00178713;
         'd3852: data <= 32'hfce42c23;         'd3853: data <= 32'hfdc42703;
         'd3854: data <= 32'h00f707b3;         'd3855: data <= 32'h03000713;
         'd3856: data <= 32'h00e78023;         'd3857: data <= 32'hfd842703;
         'd3858: data <= 32'h00042783;         'd3859: data <= 32'h02f77863;
         'd3860: data <= 32'hfd842703;         'd3861: data <= 32'h01f00793;
         'd3862: data <= 32'hfce7f8e3;         'd3863: data <= 32'h0200006f;
         'd3864: data <= 32'hfd842783;         'd3865: data <= 32'h00178713;
         'd3866: data <= 32'hfce42c23;         'd3867: data <= 32'hfdc42703;
         'd3868: data <= 32'h00f707b3;         'd3869: data <= 32'h03000713;
         'd3870: data <= 32'h00e78023;         'd3871: data <= 32'h00842783;
         'd3872: data <= 32'h0017f793;         'd3873: data <= 32'h00078e63;
         'd3874: data <= 32'hfd842703;         'd3875: data <= 32'h00442783;
         'd3876: data <= 32'h00f77863;         'd3877: data <= 32'hfd842703;
         'd3878: data <= 32'h01f00793;         'd3879: data <= 32'hfce7f2e3;
         'd3880: data <= 32'h00842783;         'd3881: data <= 32'h0107f793;
         'd3882: data <= 32'h14078063;         'd3883: data <= 32'h00842783;
         'd3884: data <= 32'h4007f793;         'd3885: data <= 32'h04079863;
         'd3886: data <= 32'hfd842783;         'd3887: data <= 32'h04078463;
         'd3888: data <= 32'hfd842703;         'd3889: data <= 32'h00042783;
         'd3890: data <= 32'h00f70863;         'd3891: data <= 32'hfd842703;
         'd3892: data <= 32'h00442783;         'd3893: data <= 32'h02f71863;
         'd3894: data <= 32'hfd842783;         'd3895: data <= 32'hfff78793;
         'd3896: data <= 32'hfcf42c23;         'd3897: data <= 32'hfd842783;
         'd3898: data <= 32'h00078e63;         'd3899: data <= 32'hfd042703;
         'd3900: data <= 32'h01000793;         'd3901: data <= 32'h00f71863;
         'd3902: data <= 32'hfd842783;         'd3903: data <= 32'hfff78793;
         'd3904: data <= 32'hfcf42c23;         'd3905: data <= 32'hfd042703;
         'd3906: data <= 32'h01000793;         'd3907: data <= 32'h02f71e63;
         'd3908: data <= 32'h00842783;         'd3909: data <= 32'h0207f793;
         'd3910: data <= 32'h02079863;         'd3911: data <= 32'hfd842703;
         'd3912: data <= 32'h01f00793;         'd3913: data <= 32'h02e7e263;
         'd3914: data <= 32'hfd842783;         'd3915: data <= 32'h00178713;
         'd3916: data <= 32'hfce42c23;         'd3917: data <= 32'hfdc42703;
         'd3918: data <= 32'h00f707b3;         'd3919: data <= 32'h07800713;
         'd3920: data <= 32'h00e78023;         'd3921: data <= 32'h07c0006f;
         'd3922: data <= 32'hfd042703;         'd3923: data <= 32'h01000793;
         'd3924: data <= 32'h02f71e63;         'd3925: data <= 32'h00842783;
         'd3926: data <= 32'h0207f793;         'd3927: data <= 32'h02078863;
         'd3928: data <= 32'hfd842703;         'd3929: data <= 32'h01f00793;
         'd3930: data <= 32'h02e7e263;         'd3931: data <= 32'hfd842783;
         'd3932: data <= 32'h00178713;         'd3933: data <= 32'hfce42c23;
         'd3934: data <= 32'hfdc42703;         'd3935: data <= 32'h00f707b3;
         'd3936: data <= 32'h05800713;         'd3937: data <= 32'h00e78023;
         'd3938: data <= 32'h0380006f;         'd3939: data <= 32'hfd042703;
         'd3940: data <= 32'h00200793;         'd3941: data <= 32'h02f71663;
         'd3942: data <= 32'hfd842703;         'd3943: data <= 32'h01f00793;
         'd3944: data <= 32'h02e7e063;         'd3945: data <= 32'hfd842783;
         'd3946: data <= 32'h00178713;         'd3947: data <= 32'hfce42c23;
         'd3948: data <= 32'hfdc42703;         'd3949: data <= 32'h00f707b3;
         'd3950: data <= 32'h06200713;         'd3951: data <= 32'h00e78023;
         'd3952: data <= 32'hfd842703;         'd3953: data <= 32'h01f00793;
         'd3954: data <= 32'h02e7e063;         'd3955: data <= 32'hfd842783;
         'd3956: data <= 32'h00178713;         'd3957: data <= 32'hfce42c23;
         'd3958: data <= 32'hfdc42703;         'd3959: data <= 32'h00f707b3;
         'd3960: data <= 32'h03000713;         'd3961: data <= 32'h00e78023;
         'd3962: data <= 32'hfd842703;         'd3963: data <= 32'h01f00793;
         'd3964: data <= 32'h08e7e063;         'd3965: data <= 32'hfd744783;
         'd3966: data <= 32'h02078263;         'd3967: data <= 32'hfd842783;
         'd3968: data <= 32'h00178713;         'd3969: data <= 32'hfce42c23;
         'd3970: data <= 32'hfdc42703;         'd3971: data <= 32'h00f707b3;
         'd3972: data <= 32'h02d00713;         'd3973: data <= 32'h00e78023;
         'd3974: data <= 32'h0580006f;         'd3975: data <= 32'h00842783;
         'd3976: data <= 32'h0047f793;         'd3977: data <= 32'h02078263;
         'd3978: data <= 32'hfd842783;         'd3979: data <= 32'h00178713;
         'd3980: data <= 32'hfce42c23;         'd3981: data <= 32'hfdc42703;
         'd3982: data <= 32'h00f707b3;         'd3983: data <= 32'h02b00713;
         'd3984: data <= 32'h00e78023;         'd3985: data <= 32'h02c0006f;
         'd3986: data <= 32'h00842783;         'd3987: data <= 32'h0087f793;
         'd3988: data <= 32'h02078063;         'd3989: data <= 32'hfd842783;
         'd3990: data <= 32'h00178713;         'd3991: data <= 32'hfce42c23;
         'd3992: data <= 32'hfdc42703;         'd3993: data <= 32'h00f707b3;
         'd3994: data <= 32'h02000713;         'd3995: data <= 32'h00e78023;
         'd3996: data <= 32'h00842883;         'd3997: data <= 32'h00442803;
         'd3998: data <= 32'hfd842783;         'd3999: data <= 32'hfdc42703;
         'd4000: data <= 32'hfe042683;         'd4001: data <= 32'hfe442603;
         'd4002: data <= 32'hfe842583;         'd4003: data <= 32'hfec42503;
         'd4004: data <= 32'hbe1ff0ef;         'd4005: data <= 32'h00050793;
         'd4006: data <= 32'h00078513;         'd4007: data <= 32'h02c12083;
         'd4008: data <= 32'h02812403;         'd4009: data <= 32'h03010113;
         'd4010: data <= 32'h00008067;         'd4011: data <= 32'hf9010113;
         'd4012: data <= 32'h06112623;         'd4013: data <= 32'h06812423;
         'd4014: data <= 32'h07010413;         'd4015: data <= 32'hfaa42e23;
         'd4016: data <= 32'hfab42c23;         'd4017: data <= 32'hfac42a23;
         'd4018: data <= 32'hfad42823;         'd4019: data <= 32'hfae42623;
         'd4020: data <= 32'hfb042223;         'd4021: data <= 32'hfb142023;
         'd4022: data <= 32'hfaf405a3;         'd4023: data <= 32'hfe042623;
         'd4024: data <= 32'hfac42783;         'd4025: data <= 32'h00079863;
         'd4026: data <= 32'h00442783;         'd4027: data <= 32'hfef7f793;
         'd4028: data <= 32'h00f42223;         'd4029: data <= 32'h00442783;
         'd4030: data <= 32'h4007f793;         'd4031: data <= 32'h00078663;
         'd4032: data <= 32'hfac42783;         'd4033: data <= 32'h0a078263;
         'd4034: data <= 32'hfac42783;         'd4035: data <= 32'hfa442583;
         'd4036: data <= 32'h00078513;         'd4037: data <= 32'h08c010ef;
         'd4038: data <= 32'h00050793;         'd4039: data <= 32'hfef405a3;
         'd4040: data <= 32'hfeb44703;         'd4041: data <= 32'h00900793;
         'd4042: data <= 32'h00e7ea63;         'd4043: data <= 32'hfeb44783;
         'd4044: data <= 32'h03078793;         'd4045: data <= 32'h0ff7f793;
         'd4046: data <= 32'h0300006f;         'd4047: data <= 32'h00442783;
         'd4048: data <= 32'h0207f793;         'd4049: data <= 32'h00078663;
         'd4050: data <= 32'h04100793;         'd4051: data <= 32'h0080006f;
         'd4052: data <= 32'h06100793;         'd4053: data <= 32'hfeb44703;
         'd4054: data <= 32'h00e787b3;         'd4055: data <= 32'h0ff7f793;
         'd4056: data <= 32'hff678793;         'd4057: data <= 32'h0ff7f793;
         'd4058: data <= 32'hfec42703;         'd4059: data <= 32'h00170693;
         'd4060: data <= 32'hfed42623;         'd4061: data <= 32'hff040693;
         'd4062: data <= 32'h00e68733;         'd4063: data <= 32'hfcf70c23;
         'd4064: data <= 32'hfa442583;         'd4065: data <= 32'hfac42503;
         'd4066: data <= 32'h7d1000ef;         'd4067: data <= 32'h00050793;
         'd4068: data <= 32'hfaf42623;         'd4069: data <= 32'hfac42783;
         'd4070: data <= 32'h00078863;         'd4071: data <= 32'hfec42703;
         'd4072: data <= 32'h01f00793;         'd4073: data <= 32'hf6e7f2e3;
         'd4074: data <= 32'hfab44683;         'd4075: data <= 32'hfc840713;
         'd4076: data <= 32'h00442783;         'd4077: data <= 32'h00f12423;
         'd4078: data <= 32'h00042783;         'd4079: data <= 32'h00f12223;
         'd4080: data <= 32'hfa042783;         'd4081: data <= 32'h00f12023;
         'd4082: data <= 32'hfa442883;         'd4083: data <= 32'h00068813;
         'd4084: data <= 32'hfec42783;         'd4085: data <= 32'hfb042683;
         'd4086: data <= 32'hfb442603;         'd4087: data <= 32'hfb842583;
         'd4088: data <= 32'hfbc42503;         'd4089: data <= 32'hbcdff0ef;
         'd4090: data <= 32'h00050793;         'd4091: data <= 32'h00078513;
         'd4092: data <= 32'h06c12083;         'd4093: data <= 32'h06812403;
         'd4094: data <= 32'h07010113;         'd4095: data <= 32'h00008067;
         'd4096: data <= 32'hf8010113;         'd4097: data <= 32'h06112e23;
         'd4098: data <= 32'h06812c23;         'd4099: data <= 32'h08010413;
         'd4100: data <= 32'hfaa42623;         'd4101: data <= 32'hfab42423;
         'd4102: data <= 32'hfac42223;         'd4103: data <= 32'hfad42023;
         'd4104: data <= 32'hf8e42e23;         'd4105: data <= 32'hfc042e23;
         'd4106: data <= 32'hfa842783;         'd4107: data <= 32'h20079ee3;
         'd4108: data <= 32'h800047b7;         'd4109: data <= 32'h85478793;
         'd4110: data <= 32'hfaf42623;         'd4111: data <= 32'h20d0006f;
         'd4112: data <= 32'hfa042783;         'd4113: data <= 32'h0007c703;
         'd4114: data <= 32'h02500793;         'd4115: data <= 32'h02f70e63;
         'd4116: data <= 32'hfa042783;         'd4117: data <= 32'h0007c503;
         'd4118: data <= 32'hfdc42783;         'd4119: data <= 32'h00178713;
         'd4120: data <= 32'hfce42e23;         'd4121: data <= 32'hfac42703;
         'd4122: data <= 32'hfa442683;         'd4123: data <= 32'h00078613;
         'd4124: data <= 32'hfa842583;         'd4125: data <= 32'h000700e7;
         'd4126: data <= 32'hfa042783;         'd4127: data <= 32'h00178793;
         'd4128: data <= 32'hfaf42023;         'd4129: data <= 32'h1c50006f;
         'd4130: data <= 32'hfa042783;         'd4131: data <= 32'h00178793;
         'd4132: data <= 32'hfaf42023;         'd4133: data <= 32'hfe042623;
         'd4134: data <= 32'hfa042783;         'd4135: data <= 32'h0007c783;
         'd4136: data <= 32'hfe078793;         'd4137: data <= 32'h01000713;
         'd4138: data <= 32'h0cf76863;         'd4139: data <= 32'h00279713;
         'd4140: data <= 32'h800057b7;         'd4141: data <= 32'h64078793;
         'd4142: data <= 32'h00f707b3;         'd4143: data <= 32'h0007a783;
         'd4144: data <= 32'h00078067;         'd4145: data <= 32'hfec42783;
         'd4146: data <= 32'h0017e793;         'd4147: data <= 32'hfef42623;
         'd4148: data <= 32'hfa042783;         'd4149: data <= 32'h00178793;
         'd4150: data <= 32'hfaf42023;         'd4151: data <= 32'h00100793;
         'd4152: data <= 32'hfef42023;         'd4153: data <= 32'h09c0006f;
         'd4154: data <= 32'hfec42783;         'd4155: data <= 32'h0027e793;
         'd4156: data <= 32'hfef42623;         'd4157: data <= 32'hfa042783;
         'd4158: data <= 32'h00178793;         'd4159: data <= 32'hfaf42023;
         'd4160: data <= 32'h00100793;         'd4161: data <= 32'hfef42023;
         'd4162: data <= 32'h0780006f;         'd4163: data <= 32'hfec42783;
         'd4164: data <= 32'h0047e793;         'd4165: data <= 32'hfef42623;
         'd4166: data <= 32'hfa042783;         'd4167: data <= 32'h00178793;
         'd4168: data <= 32'hfaf42023;         'd4169: data <= 32'h00100793;
         'd4170: data <= 32'hfef42023;         'd4171: data <= 32'h0540006f;
         'd4172: data <= 32'hfec42783;         'd4173: data <= 32'h0087e793;
         'd4174: data <= 32'hfef42623;         'd4175: data <= 32'hfa042783;
         'd4176: data <= 32'h00178793;         'd4177: data <= 32'hfaf42023;
         'd4178: data <= 32'h00100793;         'd4179: data <= 32'hfef42023;
         'd4180: data <= 32'h0300006f;         'd4181: data <= 32'hfec42783;
         'd4182: data <= 32'h0107e793;         'd4183: data <= 32'hfef42623;
         'd4184: data <= 32'hfa042783;         'd4185: data <= 32'h00178793;
         'd4186: data <= 32'hfaf42023;         'd4187: data <= 32'h00100793;
         'd4188: data <= 32'hfef42023;         'd4189: data <= 32'h00c0006f;
         'd4190: data <= 32'hfe042023;         'd4191: data <= 32'h00000013;
         'd4192: data <= 32'hfe042783;         'd4193: data <= 32'hf0079ae3;
         'd4194: data <= 32'hfe042423;         'd4195: data <= 32'hfa042783;
         'd4196: data <= 32'h0007c783;         'd4197: data <= 32'h00078513;
         'd4198: data <= 32'hffcff0ef;         'd4199: data <= 32'h00050793;
         'd4200: data <= 32'h00078c63;         'd4201: data <= 32'hfa040793;
         'd4202: data <= 32'h00078513;         'd4203: data <= 32'h839ff0ef;
         'd4204: data <= 32'hfea42423;         'd4205: data <= 32'h0600006f;
         'd4206: data <= 32'hfa042783;         'd4207: data <= 32'h0007c703;
         'd4208: data <= 32'h02a00793;         'd4209: data <= 32'h04f71863;
         'd4210: data <= 32'hf9c42783;         'd4211: data <= 32'h00478713;
         'd4212: data <= 32'hf8e42e23;         'd4213: data <= 32'h0007a783;
         'd4214: data <= 32'hfcf42423;         'd4215: data <= 32'hfc842783;
         'd4216: data <= 32'h0207d063;         'd4217: data <= 32'hfec42783;
         'd4218: data <= 32'h0027e793;         'd4219: data <= 32'hfef42623;
         'd4220: data <= 32'hfc842783;         'd4221: data <= 32'h40f007b3;
         'd4222: data <= 32'hfef42423;         'd4223: data <= 32'h00c0006f;
         'd4224: data <= 32'hfc842783;         'd4225: data <= 32'hfef42423;
         'd4226: data <= 32'hfa042783;         'd4227: data <= 32'h00178793;
         'd4228: data <= 32'hfaf42023;         'd4229: data <= 32'hfe042223;
         'd4230: data <= 32'hfa042783;         'd4231: data <= 32'h0007c703;
         'd4232: data <= 32'h02e00793;         'd4233: data <= 32'h08f71463;
         'd4234: data <= 32'hfec42783;         'd4235: data <= 32'h4007e793;
         'd4236: data <= 32'hfef42623;         'd4237: data <= 32'hfa042783;
         'd4238: data <= 32'h00178793;         'd4239: data <= 32'hfaf42023;
         'd4240: data <= 32'hfa042783;         'd4241: data <= 32'h0007c783;
         'd4242: data <= 32'h00078513;         'd4243: data <= 32'hf48ff0ef;
         'd4244: data <= 32'h00050793;         'd4245: data <= 32'h00078c63;
         'd4246: data <= 32'hfa040793;         'd4247: data <= 32'h00078513;
         'd4248: data <= 32'hf84ff0ef;         'd4249: data <= 32'hfea42223;
         'd4250: data <= 32'h0440006f;         'd4251: data <= 32'hfa042783;
         'd4252: data <= 32'h0007c703;         'd4253: data <= 32'h02a00793;
         'd4254: data <= 32'h02f71a63;         'd4255: data <= 32'hf9c42783;
         'd4256: data <= 32'h00478713;         'd4257: data <= 32'hf8e42e23;
         'd4258: data <= 32'h0007a783;         'd4259: data <= 32'hfcf42223;
         'd4260: data <= 32'hfc442783;         'd4261: data <= 32'h0007d463;
         'd4262: data <= 32'h00000793;         'd4263: data <= 32'hfef42223;
         'd4264: data <= 32'hfa042783;         'd4265: data <= 32'h00178793;
         'd4266: data <= 32'hfaf42023;         'd4267: data <= 32'hfa042783;
         'd4268: data <= 32'h0007c783;         'd4269: data <= 32'hf9878793;
         'd4270: data <= 32'h01200713;         'd4271: data <= 32'h0ef76c63;
         'd4272: data <= 32'h00279713;         'd4273: data <= 32'h800057b7;
         'd4274: data <= 32'h68478793;         'd4275: data <= 32'h00f707b3;
         'd4276: data <= 32'h0007a783;         'd4277: data <= 32'h00078067;
         'd4278: data <= 32'hfec42783;         'd4279: data <= 32'h1007e793;
         'd4280: data <= 32'hfef42623;         'd4281: data <= 32'hfa042783;
         'd4282: data <= 32'h00178793;         'd4283: data <= 32'hfaf42023;
         'd4284: data <= 32'hfa042783;         'd4285: data <= 32'h0007c703;
         'd4286: data <= 32'h06c00793;         'd4287: data <= 32'h0cf71063;
         'd4288: data <= 32'hfec42783;         'd4289: data <= 32'h2007e793;
         'd4290: data <= 32'hfef42623;         'd4291: data <= 32'hfa042783;
         'd4292: data <= 32'h00178793;         'd4293: data <= 32'hfaf42023;
         'd4294: data <= 32'h0a40006f;         'd4295: data <= 32'hfec42783;
         'd4296: data <= 32'h0807e793;         'd4297: data <= 32'hfef42623;
         'd4298: data <= 32'hfa042783;         'd4299: data <= 32'h00178793;
         'd4300: data <= 32'hfaf42023;         'd4301: data <= 32'hfa042783;
         'd4302: data <= 32'h0007c703;         'd4303: data <= 32'h06800793;
         'd4304: data <= 32'h08f71263;         'd4305: data <= 32'hfec42783;
         'd4306: data <= 32'h0407e793;         'd4307: data <= 32'hfef42623;
         'd4308: data <= 32'hfa042783;         'd4309: data <= 32'h00178793;
         'd4310: data <= 32'hfaf42023;         'd4311: data <= 32'h0680006f;
         'd4312: data <= 32'hfec42783;         'd4313: data <= 32'h1007e793;
         'd4314: data <= 32'hfef42623;         'd4315: data <= 32'hfa042783;
         'd4316: data <= 32'h00178793;         'd4317: data <= 32'hfaf42023;
         'd4318: data <= 32'h0500006f;         'd4319: data <= 32'hfec42783;
         'd4320: data <= 32'h2007e793;         'd4321: data <= 32'hfef42623;
         'd4322: data <= 32'hfa042783;         'd4323: data <= 32'h00178793;
         'd4324: data <= 32'hfaf42023;         'd4325: data <= 32'h0340006f;
         'd4326: data <= 32'hfec42783;         'd4327: data <= 32'h1007e793;
         'd4328: data <= 32'hfef42623;         'd4329: data <= 32'hfa042783;
         'd4330: data <= 32'h00178793;         'd4331: data <= 32'hfaf42023;
         'd4332: data <= 32'h0180006f;         'd4333: data <= 32'h00000013;
         'd4334: data <= 32'h0100006f;         'd4335: data <= 32'h00000013;
         'd4336: data <= 32'h0080006f;         'd4337: data <= 32'h00000013;
         'd4338: data <= 32'hfa042783;         'd4339: data <= 32'h0007c783;
         'd4340: data <= 32'hfdb78793;         'd4341: data <= 32'h05300713;
         'd4342: data <= 32'h62f76c63;         'd4343: data <= 32'h00279713;
         'd4344: data <= 32'h800057b7;         'd4345: data <= 32'h6d078793;
         'd4346: data <= 32'h00f707b3;         'd4347: data <= 32'h0007a783;
         'd4348: data <= 32'h00078067;         'd4349: data <= 32'hfa042783;
         'd4350: data <= 32'h0007c703;         'd4351: data <= 32'h07800793;
         'd4352: data <= 32'h00f70a63;         'd4353: data <= 32'hfa042783;
         'd4354: data <= 32'h0007c703;         'd4355: data <= 32'h05800793;
         'd4356: data <= 32'h00f71863;         'd4357: data <= 32'h01000793;
         'd4358: data <= 32'hfcf42c23;         'd4359: data <= 32'h0500006f;
         'd4360: data <= 32'hfa042783;         'd4361: data <= 32'h0007c703;
         'd4362: data <= 32'h06f00793;         'd4363: data <= 32'h00f71863;
         'd4364: data <= 32'h00800793;         'd4365: data <= 32'hfcf42c23;
         'd4366: data <= 32'h0340006f;         'd4367: data <= 32'hfa042783;
         'd4368: data <= 32'h0007c703;         'd4369: data <= 32'h06200793;
         'd4370: data <= 32'h00f71863;         'd4371: data <= 32'h00200793;
         'd4372: data <= 32'hfcf42c23;         'd4373: data <= 32'h0180006f;
         'd4374: data <= 32'h00a00793;         'd4375: data <= 32'hfcf42c23;
         'd4376: data <= 32'hfec42783;         'd4377: data <= 32'hfef7f793;
         'd4378: data <= 32'hfef42623;         'd4379: data <= 32'hfa042783;
         'd4380: data <= 32'h0007c703;         'd4381: data <= 32'h05800793;
         'd4382: data <= 32'h00f71863;         'd4383: data <= 32'hfec42783;
         'd4384: data <= 32'h0207e793;         'd4385: data <= 32'hfef42623;
         'd4386: data <= 32'hfa042783;         'd4387: data <= 32'h0007c703;
         'd4388: data <= 32'h06900793;         'd4389: data <= 32'h02f70063;
         'd4390: data <= 32'hfa042783;         'd4391: data <= 32'h0007c703;
         'd4392: data <= 32'h06400793;         'd4393: data <= 32'h00f70863;
         'd4394: data <= 32'hfec42783;         'd4395: data <= 32'hff37f793;
         'd4396: data <= 32'hfef42623;         'd4397: data <= 32'hfec42783;
         'd4398: data <= 32'h4007f793;         'd4399: data <= 32'h00078863;
         'd4400: data <= 32'hfec42783;         'd4401: data <= 32'hffe7f793;
         'd4402: data <= 32'hfef42623;         'd4403: data <= 32'hfa042783;
         'd4404: data <= 32'h0007c703;         'd4405: data <= 32'h06900793;
         'd4406: data <= 32'h00f70a63;         'd4407: data <= 32'hfa042783;
         'd4408: data <= 32'h0007c703;         'd4409: data <= 32'h06400793;
         'd4410: data <= 32'h14f71863;         'd4411: data <= 32'hfec42783;
         'd4412: data <= 32'h2007f793;         'd4413: data <= 32'h22079e63;
         'd4414: data <= 32'hfec42783;         'd4415: data <= 32'h1007f793;
         'd4416: data <= 32'h06078c63;         'd4417: data <= 32'hf9c42783;
         'd4418: data <= 32'h00478713;         'd4419: data <= 32'hf8e42e23;
         'd4420: data <= 32'h0007a783;         'd4421: data <= 32'hfaf42c23;
         'd4422: data <= 32'hfb842783;         'd4423: data <= 32'h41f7d713;
         'd4424: data <= 32'hfb842783;         'd4425: data <= 32'h00f747b3;
         'd4426: data <= 32'h40e787b3;         'd4427: data <= 32'h00078693;
         'd4428: data <= 32'hfb842783;         'd4429: data <= 32'h01f7d793;
         'd4430: data <= 32'h0ff7f713;         'd4431: data <= 32'hfec42783;
         'd4432: data <= 32'h00f12223;         'd4433: data <= 32'hfe842783;
         'd4434: data <= 32'h00f12023;         'd4435: data <= 32'hfe442883;
         'd4436: data <= 32'hfd842803;         'd4437: data <= 32'h00070793;
         'd4438: data <= 32'h00068713;         'd4439: data <= 32'hfa442683;
         'd4440: data <= 32'hfdc42603;         'd4441: data <= 32'hfa842583;
         'd4442: data <= 32'hfac42503;         'd4443: data <= 32'h941ff0ef;
         'd4444: data <= 32'hfca42e23;         'd4445: data <= 32'h1bc0006f;
         'd4446: data <= 32'hfec42783;         'd4447: data <= 32'h0407f793;
         'd4448: data <= 32'h00078e63;         'd4449: data <= 32'hf9c42783;
         'd4450: data <= 32'h00478713;         'd4451: data <= 32'hf8e42e23;
         'd4452: data <= 32'h0007a783;         'd4453: data <= 32'h0ff7f793;
         'd4454: data <= 32'h03c0006f;         'd4455: data <= 32'hfec42783;
         'd4456: data <= 32'h0807f793;         'd4457: data <= 32'h02078063;
         'd4458: data <= 32'hf9c42783;         'd4459: data <= 32'h00478713;
         'd4460: data <= 32'hf8e42e23;         'd4461: data <= 32'h0007a783;
         'd4462: data <= 32'h01079793;         'd4463: data <= 32'h4107d793;
         'd4464: data <= 32'h0140006f;         'd4465: data <= 32'hf9c42783;
         'd4466: data <= 32'h00478713;         'd4467: data <= 32'hf8e42e23;
         'd4468: data <= 32'h0007a783;         'd4469: data <= 32'hfaf42e23;
         'd4470: data <= 32'hfbc42783;         'd4471: data <= 32'h41f7d713;
         'd4472: data <= 32'hfbc42783;         'd4473: data <= 32'h00f747b3;
         'd4474: data <= 32'h40e787b3;         'd4475: data <= 32'h00078693;
         'd4476: data <= 32'hfbc42783;         'd4477: data <= 32'h01f7d793;
         'd4478: data <= 32'h0ff7f713;         'd4479: data <= 32'hfec42783;
         'd4480: data <= 32'h00f12223;         'd4481: data <= 32'hfe842783;
         'd4482: data <= 32'h00f12023;         'd4483: data <= 32'hfe442883;
         'd4484: data <= 32'hfd842803;         'd4485: data <= 32'h00070793;
         'd4486: data <= 32'h00068713;         'd4487: data <= 32'hfa442683;
         'd4488: data <= 32'hfdc42603;         'd4489: data <= 32'hfa842583;
         'd4490: data <= 32'hfac42503;         'd4491: data <= 32'h881ff0ef;
         'd4492: data <= 32'hfca42e23;         'd4493: data <= 32'h0fc0006f;
         'd4494: data <= 32'hfec42783;         'd4495: data <= 32'h2007f793;
         'd4496: data <= 32'h0e079863;         'd4497: data <= 32'hfec42783;
         'd4498: data <= 32'h1007f793;         'd4499: data <= 32'h04078663;
         'd4500: data <= 32'hf9c42783;         'd4501: data <= 32'h00478713;
         'd4502: data <= 32'hf8e42e23;         'd4503: data <= 32'h0007a703;
         'd4504: data <= 32'hfec42783;         'd4505: data <= 32'h00f12223;
         'd4506: data <= 32'hfe842783;         'd4507: data <= 32'h00f12023;
         'd4508: data <= 32'hfe442883;         'd4509: data <= 32'hfd842803;
         'd4510: data <= 32'h00000793;         'd4511: data <= 32'hfa442683;
         'd4512: data <= 32'hfdc42603;         'd4513: data <= 32'hfa842583;
         'd4514: data <= 32'hfac42503;         'd4515: data <= 32'h821ff0ef;
         'd4516: data <= 32'hfca42e23;         'd4517: data <= 32'h09c0006f;
         'd4518: data <= 32'hfec42783;         'd4519: data <= 32'h0407f793;
         'd4520: data <= 32'h00078e63;         'd4521: data <= 32'hf9c42783;
         'd4522: data <= 32'h00478713;         'd4523: data <= 32'hf8e42e23;
         'd4524: data <= 32'h0007a783;         'd4525: data <= 32'h0ff7f793;
         'd4526: data <= 32'h03c0006f;         'd4527: data <= 32'hfec42783;
         'd4528: data <= 32'h0807f793;         'd4529: data <= 32'h02078063;
         'd4530: data <= 32'hf9c42783;         'd4531: data <= 32'h00478713;
         'd4532: data <= 32'hf8e42e23;         'd4533: data <= 32'h0007a783;
         'd4534: data <= 32'h01079793;         'd4535: data <= 32'h0107d793;
         'd4536: data <= 32'h0140006f;         'd4537: data <= 32'hf9c42783;
         'd4538: data <= 32'h00478713;         'd4539: data <= 32'hf8e42e23;
         'd4540: data <= 32'h0007a783;         'd4541: data <= 32'hfcf42023;
         'd4542: data <= 32'hfec42783;         'd4543: data <= 32'h00f12223;
         'd4544: data <= 32'hfe842783;         'd4545: data <= 32'h00f12023;
         'd4546: data <= 32'hfe442883;         'd4547: data <= 32'hfd842803;
         'd4548: data <= 32'h00000793;         'd4549: data <= 32'hfc042703;
         'd4550: data <= 32'hfa442683;         'd4551: data <= 32'hfdc42603;
         'd4552: data <= 32'hfa842583;         'd4553: data <= 32'hfac42503;
         'd4554: data <= 32'hf84ff0ef;         'd4555: data <= 32'hfca42e23;
         'd4556: data <= 32'hfa042783;         'd4557: data <= 32'h00178793;
         'd4558: data <= 32'hfaf42023;         'd4559: data <= 32'h30c0006f;
         'd4560: data <= 32'h00100793;         'd4561: data <= 32'hfcf42a23;
         'd4562: data <= 32'hfec42783;         'd4563: data <= 32'h0027f793;
         'd4564: data <= 32'h04079063;         'd4565: data <= 32'h0280006f;
         'd4566: data <= 32'hfdc42783;         'd4567: data <= 32'h00178713;
         'd4568: data <= 32'hfce42e23;         'd4569: data <= 32'hfac42703;
         'd4570: data <= 32'hfa442683;         'd4571: data <= 32'h00078613;
         'd4572: data <= 32'hfa842583;         'd4573: data <= 32'h02000513;
         'd4574: data <= 32'h000700e7;         'd4575: data <= 32'hfd442783;
         'd4576: data <= 32'h00178713;         'd4577: data <= 32'hfce42a23;
         'd4578: data <= 32'hfe842703;         'd4579: data <= 32'hfce7e6e3;
         'd4580: data <= 32'hf9c42783;         'd4581: data <= 32'h00478713;
         'd4582: data <= 32'hf8e42e23;         'd4583: data <= 32'h0007a783;
         'd4584: data <= 32'h0ff7f513;         'd4585: data <= 32'hfdc42783;
         'd4586: data <= 32'h00178713;         'd4587: data <= 32'hfce42e23;
         'd4588: data <= 32'hfac42703;         'd4589: data <= 32'hfa442683;
         'd4590: data <= 32'h00078613;         'd4591: data <= 32'hfa842583;
         'd4592: data <= 32'h000700e7;         'd4593: data <= 32'hfec42783;
         'd4594: data <= 32'h0027f793;         'd4595: data <= 32'h04078063;
         'd4596: data <= 32'h0280006f;         'd4597: data <= 32'hfdc42783;
         'd4598: data <= 32'h00178713;         'd4599: data <= 32'hfce42e23;
         'd4600: data <= 32'hfac42703;         'd4601: data <= 32'hfa442683;
         'd4602: data <= 32'h00078613;         'd4603: data <= 32'hfa842583;
         'd4604: data <= 32'h02000513;         'd4605: data <= 32'h000700e7;
         'd4606: data <= 32'hfd442783;         'd4607: data <= 32'h00178713;
         'd4608: data <= 32'hfce42a23;         'd4609: data <= 32'hfe842703;
         'd4610: data <= 32'hfce7e6e3;         'd4611: data <= 32'hfa042783;
         'd4612: data <= 32'h00178793;         'd4613: data <= 32'hfaf42023;
         'd4614: data <= 32'h2300006f;         'd4615: data <= 32'hf9c42783;
         'd4616: data <= 32'h00478713;         'd4617: data <= 32'hf8e42e23;
         'd4618: data <= 32'h0007a783;         'd4619: data <= 32'hfcf42823;
         'd4620: data <= 32'hfe442783;         'd4621: data <= 32'h00078663;
         'd4622: data <= 32'hfe442783;         'd4623: data <= 32'h0080006f;
         'd4624: data <= 32'hfff00793;         'd4625: data <= 32'h00078593;
         'd4626: data <= 32'hfd042503;         'd4627: data <= 32'h8e4ff0ef;
         'd4628: data <= 32'hfca42623;         'd4629: data <= 32'hfec42783;
         'd4630: data <= 32'h4007f793;         'd4631: data <= 32'h00078c63;
         'd4632: data <= 32'hfcc42703;         'd4633: data <= 32'hfe442783;
         'd4634: data <= 32'h00f77463;         'd4635: data <= 32'h00070793;
         'd4636: data <= 32'hfcf42623;         'd4637: data <= 32'hfec42783;
         'd4638: data <= 32'h0027f793;         'd4639: data <= 32'h06079a63;
         'd4640: data <= 32'h0280006f;         'd4641: data <= 32'hfdc42783;
         'd4642: data <= 32'h00178713;         'd4643: data <= 32'hfce42e23;
         'd4644: data <= 32'hfac42703;         'd4645: data <= 32'hfa442683;
         'd4646: data <= 32'h00078613;         'd4647: data <= 32'hfa842583;
         'd4648: data <= 32'h02000513;         'd4649: data <= 32'h000700e7;
         'd4650: data <= 32'hfcc42783;         'd4651: data <= 32'h00178713;
         'd4652: data <= 32'hfce42623;         'd4653: data <= 32'hfe842703;
         'd4654: data <= 32'hfce7e6e3;         'd4655: data <= 32'h0340006f;
         'd4656: data <= 32'hfd042783;         'd4657: data <= 32'h00178713;
         'd4658: data <= 32'hfce42823;         'd4659: data <= 32'h0007c503;
         'd4660: data <= 32'hfdc42783;         'd4661: data <= 32'h00178713;
         'd4662: data <= 32'hfce42e23;         'd4663: data <= 32'hfac42703;
         'd4664: data <= 32'hfa442683;         'd4665: data <= 32'h00078613;
         'd4666: data <= 32'hfa842583;         'd4667: data <= 32'h000700e7;
         'd4668: data <= 32'hfd042783;         'd4669: data <= 32'h0007c783;
         'd4670: data <= 32'h02078063;         'd4671: data <= 32'hfec42783;
         'd4672: data <= 32'h4007f793;         'd4673: data <= 32'hfa078ee3;
         'd4674: data <= 32'hfe442783;         'd4675: data <= 32'hfff78713;
         'd4676: data <= 32'hfee42223;         'd4677: data <= 32'hfa0796e3;
         'd4678: data <= 32'hfec42783;         'd4679: data <= 32'h0027f793;
         'd4680: data <= 32'h04078063;         'd4681: data <= 32'h0280006f;
         'd4682: data <= 32'hfdc42783;         'd4683: data <= 32'h00178713;
         'd4684: data <= 32'hfce42e23;         'd4685: data <= 32'hfac42703;
         'd4686: data <= 32'hfa442683;         'd4687: data <= 32'h00078613;
         'd4688: data <= 32'hfa842583;         'd4689: data <= 32'h02000513;
         'd4690: data <= 32'h000700e7;         'd4691: data <= 32'hfcc42783;
         'd4692: data <= 32'h00178713;         'd4693: data <= 32'hfce42623;
         'd4694: data <= 32'hfe842703;         'd4695: data <= 32'hfce7e6e3;
         'd4696: data <= 32'hfa042783;         'd4697: data <= 32'h00178793;
         'd4698: data <= 32'hfaf42023;         'd4699: data <= 32'h0dc0006f;
         'd4700: data <= 32'h00800793;         'd4701: data <= 32'hfef42423;
         'd4702: data <= 32'hfec42783;         'd4703: data <= 32'h0217e793;
         'd4704: data <= 32'hfef42623;         'd4705: data <= 32'hf9c42783;
         'd4706: data <= 32'h00478713;         'd4707: data <= 32'hf8e42e23;
         'd4708: data <= 32'h0007a783;         'd4709: data <= 32'h00078713;
         'd4710: data <= 32'hfec42783;         'd4711: data <= 32'h00f12223;
         'd4712: data <= 32'hfe842783;         'd4713: data <= 32'h00f12023;
         'd4714: data <= 32'hfe442883;         'd4715: data <= 32'h01000813;
         'd4716: data <= 32'h00000793;         'd4717: data <= 32'hfa442683;
         'd4718: data <= 32'hfdc42603;         'd4719: data <= 32'hfa842583;
         'd4720: data <= 32'hfac42503;         'd4721: data <= 32'hce8ff0ef;
         'd4722: data <= 32'hfca42e23;         'd4723: data <= 32'hfa042783;
         'd4724: data <= 32'h00178793;         'd4725: data <= 32'hfaf42023;
         'd4726: data <= 32'h0700006f;         'd4727: data <= 32'hfdc42783;
         'd4728: data <= 32'h00178713;         'd4729: data <= 32'hfce42e23;
         'd4730: data <= 32'hfac42703;         'd4731: data <= 32'hfa442683;
         'd4732: data <= 32'h00078613;         'd4733: data <= 32'hfa842583;
         'd4734: data <= 32'h02500513;         'd4735: data <= 32'h000700e7;
         'd4736: data <= 32'hfa042783;         'd4737: data <= 32'h00178793;
         'd4738: data <= 32'hfaf42023;         'd4739: data <= 32'h03c0006f;
         'd4740: data <= 32'hfa042783;         'd4741: data <= 32'h0007c503;
         'd4742: data <= 32'hfdc42783;         'd4743: data <= 32'h00178713;
         'd4744: data <= 32'hfce42e23;         'd4745: data <= 32'hfac42703;
         'd4746: data <= 32'hfa442683;         'd4747: data <= 32'h00078613;
         'd4748: data <= 32'hfa842583;         'd4749: data <= 32'h000700e7;
         'd4750: data <= 32'hfa042783;         'd4751: data <= 32'h00178793;
         'd4752: data <= 32'hfaf42023;         'd4753: data <= 32'h00000013;
         'd4754: data <= 32'hfa042783;         'd4755: data <= 32'h0007c783;
         'd4756: data <= 32'hde079863;         'd4757: data <= 32'hfdc42703;
         'd4758: data <= 32'hfa442783;         'd4759: data <= 32'h00f76863;
         'd4760: data <= 32'hfa442783;         'd4761: data <= 32'hfff78793;
         'd4762: data <= 32'h0080006f;         'd4763: data <= 32'hfdc42783;
         'd4764: data <= 32'hfac42703;         'd4765: data <= 32'hfa442683;
         'd4766: data <= 32'h00078613;         'd4767: data <= 32'hfa842583;
         'd4768: data <= 32'h00000513;         'd4769: data <= 32'h000700e7;
         'd4770: data <= 32'hfdc42783;         'd4771: data <= 32'h00078513;
         'd4772: data <= 32'h07c12083;         'd4773: data <= 32'h07812403;
         'd4774: data <= 32'h08010113;         'd4775: data <= 32'h00008067;
         'd4776: data <= 32'hfb010113;         'd4777: data <= 32'h02112623;
         'd4778: data <= 32'h02812423;         'd4779: data <= 32'h03010413;
         'd4780: data <= 32'hfca42e23;         'd4781: data <= 32'h00b42223;
         'd4782: data <= 32'h00c42423;         'd4783: data <= 32'h00d42623;
         'd4784: data <= 32'h00e42823;         'd4785: data <= 32'h00f42a23;
         'd4786: data <= 32'h01042c23;         'd4787: data <= 32'h01142e23;
         'd4788: data <= 32'h02040793;         'd4789: data <= 32'hfcf42c23;
         'd4790: data <= 32'hfd842783;         'd4791: data <= 32'hfe478793;
         'd4792: data <= 32'hfef42423;         'd4793: data <= 32'hfe842703;
         'd4794: data <= 32'hfe440793;         'd4795: data <= 32'hfdc42683;
         'd4796: data <= 32'hfff00613;         'd4797: data <= 32'h00078593;
         'd4798: data <= 32'h800047b7;         'd4799: data <= 32'h88478513;
         'd4800: data <= 32'hd00ff0ef;         'd4801: data <= 32'hfea42623;
         'd4802: data <= 32'hfec42783;         'd4803: data <= 32'h00078513;
         'd4804: data <= 32'h02c12083;         'd4805: data <= 32'h02812403;
         'd4806: data <= 32'h05010113;         'd4807: data <= 32'h00008067;
         'd4808: data <= 32'hfb010113;         'd4809: data <= 32'h02112623;
         'd4810: data <= 32'h02812423;         'd4811: data <= 32'h03010413;
         'd4812: data <= 32'hfca42e23;         'd4813: data <= 32'hfcb42c23;
         'd4814: data <= 32'h00c42423;         'd4815: data <= 32'h00d42623;
         'd4816: data <= 32'h00e42823;         'd4817: data <= 32'h00f42a23;
         'd4818: data <= 32'h01042c23;         'd4819: data <= 32'h01142e23;
         'd4820: data <= 32'h02040793;         'd4821: data <= 32'hfcf42a23;
         'd4822: data <= 32'hfd442783;         'd4823: data <= 32'hfe878793;
         'd4824: data <= 32'hfef42423;         'd4825: data <= 32'hfe842783;
         'd4826: data <= 32'h00078713;         'd4827: data <= 32'hfd842683;
         'd4828: data <= 32'hfff00613;         'd4829: data <= 32'hfdc42583;
         'd4830: data <= 32'h800047b7;         'd4831: data <= 32'h80478513;
         'd4832: data <= 32'hc80ff0ef;         'd4833: data <= 32'hfea42623;
         'd4834: data <= 32'hfec42783;         'd4835: data <= 32'h00078513;
         'd4836: data <= 32'h02c12083;         'd4837: data <= 32'h02812403;
         'd4838: data <= 32'h05010113;         'd4839: data <= 32'h00008067;
         'd4840: data <= 32'hfb010113;         'd4841: data <= 32'h02112623;
         'd4842: data <= 32'h02812423;         'd4843: data <= 32'h03010413;
         'd4844: data <= 32'hfca42e23;         'd4845: data <= 32'hfcb42c23;
         'd4846: data <= 32'hfcc42a23;         'd4847: data <= 32'h00d42623;
         'd4848: data <= 32'h00e42823;         'd4849: data <= 32'h00f42a23;
         'd4850: data <= 32'h01042c23;         'd4851: data <= 32'h01142e23;
         'd4852: data <= 32'h02040793;         'd4853: data <= 32'hfcf42823;
         'd4854: data <= 32'hfd042783;         'd4855: data <= 32'hfec78793;
         'd4856: data <= 32'hfef42423;         'd4857: data <= 32'hfe842783;
         'd4858: data <= 32'h00078713;         'd4859: data <= 32'hfd442683;
         'd4860: data <= 32'hfd842603;         'd4861: data <= 32'hfdc42583;
         'd4862: data <= 32'h800047b7;         'd4863: data <= 32'h80478513;
         'd4864: data <= 32'hc00ff0ef;         'd4865: data <= 32'hfea42623;
         'd4866: data <= 32'hfec42783;         'd4867: data <= 32'h00078513;
         'd4868: data <= 32'h02c12083;         'd4869: data <= 32'h02812403;
         'd4870: data <= 32'h05010113;         'd4871: data <= 32'h00008067;
         'd4872: data <= 32'hfd010113;         'd4873: data <= 32'h02112623;
         'd4874: data <= 32'h02812423;         'd4875: data <= 32'h03010413;
         'd4876: data <= 32'hfca42e23;         'd4877: data <= 32'hfcb42c23;
         'd4878: data <= 32'hfec40793;         'd4879: data <= 32'hfd842703;
         'd4880: data <= 32'hfdc42683;         'd4881: data <= 32'hfff00613;
         'd4882: data <= 32'h00078593;         'd4883: data <= 32'h800047b7;
         'd4884: data <= 32'h88478513;         'd4885: data <= 32'hbacff0ef;
         'd4886: data <= 32'h00050793;         'd4887: data <= 32'h00078513;
         'd4888: data <= 32'h02c12083;         'd4889: data <= 32'h02812403;
         'd4890: data <= 32'h03010113;         'd4891: data <= 32'h00008067;
         'd4892: data <= 32'hfe010113;         'd4893: data <= 32'h00112e23;
         'd4894: data <= 32'h00812c23;         'd4895: data <= 32'h02010413;
         'd4896: data <= 32'hfea42623;         'd4897: data <= 32'hfeb42423;
         'd4898: data <= 32'hfec42223;         'd4899: data <= 32'hfed42023;
         'd4900: data <= 32'hfe042703;         'd4901: data <= 32'hfe442683;
         'd4902: data <= 32'hfe842603;         'd4903: data <= 32'hfec42583;
         'd4904: data <= 32'h800047b7;         'd4905: data <= 32'h80478513;
         'd4906: data <= 32'hb58ff0ef;         'd4907: data <= 32'h00050793;
         'd4908: data <= 32'h00078513;         'd4909: data <= 32'h01c12083;
         'd4910: data <= 32'h01812403;         'd4911: data <= 32'h02010113;
         'd4912: data <= 32'h00008067;         'd4913: data <= 32'hfb010113;
         'd4914: data <= 32'h02112623;         'd4915: data <= 32'h02812423;
         'd4916: data <= 32'h03010413;         'd4917: data <= 32'hfca42e23;
         'd4918: data <= 32'hfcb42c23;         'd4919: data <= 32'hfcc42a23;
         'd4920: data <= 32'h00d42623;         'd4921: data <= 32'h00e42823;
         'd4922: data <= 32'h00f42a23;         'd4923: data <= 32'h01042c23;
         'd4924: data <= 32'h01142e23;         'd4925: data <= 32'h02040793;
         'd4926: data <= 32'hfcf42823;         'd4927: data <= 32'hfd042783;
         'd4928: data <= 32'hfec78793;         'd4929: data <= 32'hfef42423;
         'd4930: data <= 32'hfdc42783;         'd4931: data <= 32'hfef42023;
         'd4932: data <= 32'hfd842783;         'd4933: data <= 32'hfef42223;
         'd4934: data <= 32'hfe842703;         'd4935: data <= 32'hfe040793;
         'd4936: data <= 32'hfd442683;         'd4937: data <= 32'hfff00613;
         'd4938: data <= 32'h00078593;         'd4939: data <= 32'h800047b7;
         'd4940: data <= 32'h8d078513;         'd4941: data <= 32'haccff0ef;
         'd4942: data <= 32'hfea42623;         'd4943: data <= 32'hfec42783;
         'd4944: data <= 32'h00078513;         'd4945: data <= 32'h02c12083;
         'd4946: data <= 32'h02812403;         'd4947: data <= 32'h05010113;
         'd4948: data <= 32'h00008067;         'd4949: data <= 32'hfe010113;
         'd4950: data <= 32'h00812e23;         'd4951: data <= 32'h02010413;
         'd4952: data <= 32'h00050793;         'd4953: data <= 32'hfef407a3;
         'd4954: data <= 32'h00000013;         'd4955: data <= 32'hb00007b7;
         'd4956: data <= 32'h00478793;         'd4957: data <= 32'h0007a703;
         'd4958: data <= 32'h000107b7;         'd4959: data <= 32'h00f777b3;
         'd4960: data <= 32'hfe0786e3;         'd4961: data <= 32'hb00007b7;
         'd4962: data <= 32'h00c78793;         'd4963: data <= 32'hfef44703;
         'd4964: data <= 32'h00e7a023;         'd4965: data <= 32'h00000013;
         'd4966: data <= 32'h01c12403;         'd4967: data <= 32'h02010113;
         'd4968: data <= 32'h00008067;         'd4969: data <= 32'hfe010113;
         'd4970: data <= 32'h00812e23;         'd4971: data <= 32'h02010413;
         'd4972: data <= 32'hc00022f3;         'd4973: data <= 32'hfe542623;
         'd4974: data <= 32'h00028793;         'd4975: data <= 32'h00078513;
         'd4976: data <= 32'h01c12403;         'd4977: data <= 32'h02010113;
         'd4978: data <= 32'h00008067;         'd4979: data <= 32'hff010113;
         'd4980: data <= 32'h00112623;         'd4981: data <= 32'h00812423;
         'd4982: data <= 32'h01010413;         'd4983: data <= 32'hfc9ff0ef;
         'd4984: data <= 32'h00050713;         'd4985: data <= 32'h86e1ac23;
         'd4986: data <= 32'h00000013;         'd4987: data <= 32'h00c12083;
         'd4988: data <= 32'h00812403;         'd4989: data <= 32'h01010113;
         'd4990: data <= 32'h00008067;         'd4991: data <= 32'hff010113;
         'd4992: data <= 32'h00112623;         'd4993: data <= 32'h00812423;
         'd4994: data <= 32'h01010413;         'd4995: data <= 32'hf99ff0ef;
         'd4996: data <= 32'h00050713;         'd4997: data <= 32'h86e1ae23;
         'd4998: data <= 32'h00000013;         'd4999: data <= 32'h00c12083;
         'd5000: data <= 32'h00812403;         'd5001: data <= 32'h01010113;
         'd5002: data <= 32'h00008067;         'd5003: data <= 32'hfe010113;
         'd5004: data <= 32'h00812e23;         'd5005: data <= 32'h02010413;
         'd5006: data <= 32'h87c1a703;         'd5007: data <= 32'h8781a783;
         'd5008: data <= 32'h40f707b3;         'd5009: data <= 32'hfef42623;
         'd5010: data <= 32'hfec42783;         'd5011: data <= 32'h00078513;
         'd5012: data <= 32'h01c12403;         'd5013: data <= 32'h02010113;
         'd5014: data <= 32'h00008067;         'd5015: data <= 32'hfd010113;
         'd5016: data <= 32'h02112623;         'd5017: data <= 32'h02812423;
         'd5018: data <= 32'h03010413;         'd5019: data <= 32'hfca42e23;
         'd5020: data <= 32'hfdc42703;         'd5021: data <= 32'h02faf7b7;
         'd5022: data <= 32'h08078593;         'd5023: data <= 32'h00070513;
         'd5024: data <= 32'h0d8000ef;         'd5025: data <= 32'h00050793;
         'd5026: data <= 32'hfef42623;         'd5027: data <= 32'hfec42783;
         'd5028: data <= 32'h00078513;         'd5029: data <= 32'h02c12083;
         'd5030: data <= 32'h02812403;         'd5031: data <= 32'h03010113;
         'd5032: data <= 32'h00008067;         'd5033: data <= 32'hfe010113;
         'd5034: data <= 32'h00112e23;         'd5035: data <= 32'h00812c23;
         'd5036: data <= 32'h02010413;         'd5037: data <= 32'hfea42623;
         'd5038: data <= 32'hfeb42423;         'd5039: data <= 32'hfec42223;
         'd5040: data <= 32'hb00007b7;         'd5041: data <= 32'h1b200713;
         'd5042: data <= 32'h00e7a023;         'd5043: data <= 32'h800067b7;
         'd5044: data <= 32'h82078513;         'd5045: data <= 32'hbcdff0ef;
         'd5046: data <= 32'h800067b7;         'd5047: data <= 32'h83078513;
         'd5048: data <= 32'hbc1ff0ef;         'd5049: data <= 32'h800067b7;
         'd5050: data <= 32'h82078513;         'd5051: data <= 32'hbb5ff0ef;
         'd5052: data <= 32'hfec42783;         'd5053: data <= 32'h00100713;
         'd5054: data <= 32'h00e78023;         'd5055: data <= 32'h00000013;
         'd5056: data <= 32'h01c12083;         'd5057: data <= 32'h01812403;
         'd5058: data <= 32'h02010113;         'd5059: data <= 32'h00008067;
         'd5060: data <= 32'hfe010113;         'd5061: data <= 32'h00812e23;
         'd5062: data <= 32'h02010413;         'd5063: data <= 32'hfea42623;
         'd5064: data <= 32'hfec42783;         'd5065: data <= 32'h00078023;
         'd5066: data <= 32'h0000006f;         'd5067: data <= 32'h00050613;
         'd5068: data <= 32'h00000513;         'd5069: data <= 32'h0015f693;
         'd5070: data <= 32'h00068463;         'd5071: data <= 32'h00c50533;
         'd5072: data <= 32'h0015d593;         'd5073: data <= 32'h00161613;
         'd5074: data <= 32'hfe0596e3;         'd5075: data <= 32'h00008067;
         'd5076: data <= 32'h06054063;         'd5077: data <= 32'h0605c663;
         'd5078: data <= 32'h00058613;         'd5079: data <= 32'h00050593;
         'd5080: data <= 32'hfff00513;         'd5081: data <= 32'h02060c63;
         'd5082: data <= 32'h00100693;         'd5083: data <= 32'h00b67a63;
         'd5084: data <= 32'h00c05863;         'd5085: data <= 32'h00161613;
         'd5086: data <= 32'h00169693;         'd5087: data <= 32'hfeb66ae3;
         'd5088: data <= 32'h00000513;         'd5089: data <= 32'h00c5e663;
         'd5090: data <= 32'h40c585b3;         'd5091: data <= 32'h00d56533;
         'd5092: data <= 32'h0016d693;         'd5093: data <= 32'h00165613;
         'd5094: data <= 32'hfe0696e3;         'd5095: data <= 32'h00008067;
         'd5096: data <= 32'h00008293;         'd5097: data <= 32'hfb5ff0ef;
         'd5098: data <= 32'h00058513;         'd5099: data <= 32'h00028067;
         'd5100: data <= 32'h40a00533;         'd5101: data <= 32'h00b04863;
         'd5102: data <= 32'h40b005b3;         'd5103: data <= 32'hf9dff06f;
         'd5104: data <= 32'h40b005b3;         'd5105: data <= 32'h00008293;
         'd5106: data <= 32'hf91ff0ef;         'd5107: data <= 32'h40a00533;
         'd5108: data <= 32'h00028067;         'd5109: data <= 32'h00008293;
         'd5110: data <= 32'h0005ca63;         'd5111: data <= 32'h00054c63;
         'd5112: data <= 32'hf79ff0ef;         'd5113: data <= 32'h00058513;
         'd5114: data <= 32'h00028067;         'd5115: data <= 32'h40b005b3;
         'd5116: data <= 32'hfe0558e3;         'd5117: data <= 32'h40a00533;
         'd5118: data <= 32'hf61ff0ef;         'd5119: data <= 32'h40b00533;
         'd5120: data <= 32'h00028067;         'd5121: data <= 32'h74617453;
         'd5122: data <= 32'h00006369;         'd5123: data <= 32'h70616548;
         'd5124: data <= 32'h00000000;         'd5125: data <= 32'h63617453;
         'd5126: data <= 32'h0000006b;         'd5127: data <= 32'h70206b36;
         'd5128: data <= 32'h6f667265;         'd5129: data <= 32'h6e616d72;
         'd5130: data <= 32'h72206563;         'd5131: data <= 32'h70206e75;
         'd5132: data <= 32'h6d617261;         'd5133: data <= 32'h72657465;
         'd5134: data <= 32'h6f662073;         'd5135: data <= 32'h6f632072;
         'd5136: data <= 32'h616d6572;         'd5137: data <= 32'h0a2e6b72;
         'd5138: data <= 32'h00000000;         'd5139: data <= 32'h76206b36;
         'd5140: data <= 32'h64696c61;         'd5141: data <= 32'h6f697461;
         'd5142: data <= 32'h7572206e;         'd5143: data <= 32'h6170206e;
         'd5144: data <= 32'h656d6172;         'd5145: data <= 32'h73726574;
         'd5146: data <= 32'h726f6620;         'd5147: data <= 32'h726f6320;
         'd5148: data <= 32'h72616d65;         'd5149: data <= 32'h000a2e6b;
         'd5150: data <= 32'h666f7250;         'd5151: data <= 32'h20656c69;
         'd5152: data <= 32'h656e6567;         'd5153: data <= 32'h69746172;
         'd5154: data <= 32'h72206e6f;         'd5155: data <= 32'h70206e75;
         'd5156: data <= 32'h6d617261;         'd5157: data <= 32'h72657465;
         'd5158: data <= 32'h6f662073;         'd5159: data <= 32'h6f632072;
         'd5160: data <= 32'h616d6572;         'd5161: data <= 32'h0a2e6b72;
         'd5162: data <= 32'h00000000;         'd5163: data <= 32'h70204b32;
         'd5164: data <= 32'h6f667265;         'd5165: data <= 32'h6e616d72;
         'd5166: data <= 32'h72206563;         'd5167: data <= 32'h70206e75;
         'd5168: data <= 32'h6d617261;         'd5169: data <= 32'h72657465;
         'd5170: data <= 32'h6f662073;         'd5171: data <= 32'h6f632072;
         'd5172: data <= 32'h616d6572;         'd5173: data <= 32'h0a2e6b72;
         'd5174: data <= 32'h00000000;         'd5175: data <= 32'h76204b32;
         'd5176: data <= 32'h64696c61;         'd5177: data <= 32'h6f697461;
         'd5178: data <= 32'h7572206e;         'd5179: data <= 32'h6170206e;
         'd5180: data <= 32'h656d6172;         'd5181: data <= 32'h73726574;
         'd5182: data <= 32'h726f6620;         'd5183: data <= 32'h726f6320;
         'd5184: data <= 32'h72616d65;         'd5185: data <= 32'h000a2e6b;
         'd5186: data <= 32'h5d75255b;         'd5187: data <= 32'h4f525245;
         'd5188: data <= 32'h6c202152;         'd5189: data <= 32'h20747369;
         'd5190: data <= 32'h20637263;         'd5191: data <= 32'h30257830;
         'd5192: data <= 32'h2d207834;         'd5193: data <= 32'h6f687320;
         'd5194: data <= 32'h20646c75;         'd5195: data <= 32'h30206562;
         'd5196: data <= 32'h34302578;         'd5197: data <= 32'h00000a78;
         'd5198: data <= 32'h5d75255b;         'd5199: data <= 32'h4f525245;
         'd5200: data <= 32'h6d202152;         'd5201: data <= 32'h69727461;
         'd5202: data <= 32'h72632078;         'd5203: data <= 32'h78302063;
         'd5204: data <= 32'h78343025;         'd5205: data <= 32'h73202d20;
         'd5206: data <= 32'h6c756f68;         'd5207: data <= 32'h65622064;
         'd5208: data <= 32'h25783020;         'd5209: data <= 32'h0a783430;
         'd5210: data <= 32'h00000000;         'd5211: data <= 32'h5d75255b;
         'd5212: data <= 32'h4f525245;         'd5213: data <= 32'h73202152;
         'd5214: data <= 32'h65746174;         'd5215: data <= 32'h63726320;
         'd5216: data <= 32'h25783020;         'd5217: data <= 32'h20783430;
         'd5218: data <= 32'h6873202d;         'd5219: data <= 32'h646c756f;
         'd5220: data <= 32'h20656220;         'd5221: data <= 32'h30257830;
         'd5222: data <= 32'h000a7834;         'd5223: data <= 32'h65726f43;
         'd5224: data <= 32'h6b72614d;         'd5225: data <= 32'h7a695320;
         'd5226: data <= 32'h20202065;         'd5227: data <= 32'h25203a20;
         'd5228: data <= 32'h000a756c;         'd5229: data <= 32'h61746f54;
         'd5230: data <= 32'h6974206c;         'd5231: data <= 32'h20736b63;
         'd5232: data <= 32'h20202020;         'd5233: data <= 32'h25203a20;
         'd5234: data <= 32'h000a756c;         'd5235: data <= 32'h61746f54;
         'd5236: data <= 32'h6974206c;         'd5237: data <= 32'h2820656d;
         'd5238: data <= 32'h73636573;         'd5239: data <= 32'h25203a29;
         'd5240: data <= 32'h00000a64;         'd5241: data <= 32'h72657449;
         'd5242: data <= 32'h6f697461;         'd5243: data <= 32'h532f736e;
         'd5244: data <= 32'h20206365;         'd5245: data <= 32'h25203a20;
         'd5246: data <= 32'h00000a64;         'd5247: data <= 32'h4f525245;
         'd5248: data <= 32'h4d202152;         'd5249: data <= 32'h20747375;
         'd5250: data <= 32'h63657865;         'd5251: data <= 32'h20657475;
         'd5252: data <= 32'h20726f66;         'd5253: data <= 32'h6c207461;
         'd5254: data <= 32'h74736165;         'd5255: data <= 32'h20303120;
         'd5256: data <= 32'h73636573;         'd5257: data <= 32'h726f6620;
         'd5258: data <= 32'h76206120;         'd5259: data <= 32'h64696c61;
         'd5260: data <= 32'h73657220;         'd5261: data <= 32'h21746c75;
         'd5262: data <= 32'h0000000a;         'd5263: data <= 32'h72657449;
         'd5264: data <= 32'h6f697461;         'd5265: data <= 32'h2020736e;
         'd5266: data <= 32'h20202020;         'd5267: data <= 32'h25203a20;
         'd5268: data <= 32'h000a756c;         'd5269: data <= 32'h63736972;
         'd5270: data <= 32'h6f6e2d76;         'd5271: data <= 32'h652d656e;
         'd5272: data <= 32'h6465626d;         'd5273: data <= 32'h6363672d;
         'd5274: data <= 32'h50782820;         'd5275: data <= 32'h206b6361;
         'd5276: data <= 32'h20554e47;         'd5277: data <= 32'h43534952;
         'd5278: data <= 32'h4520562d;         'd5279: data <= 32'h6465626d;
         'd5280: data <= 32'h20646564;         'd5281: data <= 32'h20434347;
         'd5282: data <= 32'h5f363878;         'd5283: data <= 32'h20293436;
         'd5284: data <= 32'h322e3031;         'd5285: data <= 32'h0000302e;
         'd5286: data <= 32'h706d6f43;         'd5287: data <= 32'h72656c69;
         'd5288: data <= 32'h72657620;         'd5289: data <= 32'h6e6f6973;
         'd5290: data <= 32'h25203a20;         'd5291: data <= 32'h00000a73;
         'd5292: data <= 32'h20304f2d;         'd5293: data <= 32'h2d20672d;
         'd5294: data <= 32'h6372616d;         'd5295: data <= 32'h76723d68;
         'd5296: data <= 32'h20693233;         'd5297: data <= 32'h62616d2d;
         'd5298: data <= 32'h6c693d69;         'd5299: data <= 32'h20323370;
         'd5300: data <= 32'h6c61572d;         'd5301: data <= 32'h572d206c;
         'd5302: data <= 32'h752d6f6e;         'd5303: data <= 32'h6573756e;
         'd5304: data <= 32'h662d2064;         'd5305: data <= 32'h65657266;
         'd5306: data <= 32'h6e617473;         'd5307: data <= 32'h676e6964;
         'd5308: data <= 32'h732d2d20;         'd5309: data <= 32'h73636570;
         'd5310: data <= 32'h6e616e3d;         'd5311: data <= 32'h70732e6f;
         'd5312: data <= 32'h20736365;         'd5313: data <= 32'h5250442d;
         'd5314: data <= 32'h46544e49;         'd5315: data <= 32'h5349445f;
         'd5316: data <= 32'h454c4241;         'd5317: data <= 32'h5055535f;
         'd5318: data <= 32'h54524f50;         'd5319: data <= 32'h4f4c465f;
         'd5320: data <= 32'h2d205441;         'd5321: data <= 32'h49525044;
         'd5322: data <= 32'h5f46544e;         'd5323: data <= 32'h41534944;
         'd5324: data <= 32'h5f454c42;         'd5325: data <= 32'h50505553;
         'd5326: data <= 32'h5f54524f;         'd5327: data <= 32'h4f505845;
         'd5328: data <= 32'h544e454e;         'd5329: data <= 32'h204c4149;
         'd5330: data <= 32'h5250442d;         'd5331: data <= 32'h46544e49;
         'd5332: data <= 32'h5349445f;         'd5333: data <= 32'h454c4241;
         'd5334: data <= 32'h5055535f;         'd5335: data <= 32'h54524f50;
         'd5336: data <= 32'h4e4f4c5f;         'd5337: data <= 32'h4f4c5f47;
         'd5338: data <= 32'h2d20474e;         'd5339: data <= 32'h6c6c6157;
         'd5340: data <= 32'h6e572d20;         'd5341: data <= 32'h616d2d6f;
         'd5342: data <= 32'h2d206e69;         'd5343: data <= 32'h52455044;
         'd5344: data <= 32'h4d524f46;         'd5345: data <= 32'h45434e41;
         'd5346: data <= 32'h4e55525f;         'd5347: data <= 32'h2020313d;
         'd5348: data <= 32'h20304f2d;         'd5349: data <= 32'h0000672d;
         'd5350: data <= 32'h706d6f43;         'd5351: data <= 32'h72656c69;
         'd5352: data <= 32'h616c6620;         'd5353: data <= 32'h20207367;
         'd5354: data <= 32'h25203a20;         'd5355: data <= 32'h00000a73;
         'd5356: data <= 32'h43415453;         'd5357: data <= 32'h0000004b;
         'd5358: data <= 32'h6f6d654d;         'd5359: data <= 32'h6c207972;
         'd5360: data <= 32'h7461636f;         'd5361: data <= 32'h206e6f69;
         'd5362: data <= 32'h25203a20;         'd5363: data <= 32'h00000a73;
         'd5364: data <= 32'h64656573;         'd5365: data <= 32'h20637263;
         'd5366: data <= 32'h20202020;         'd5367: data <= 32'h20202020;
         'd5368: data <= 32'h30203a20;         'd5369: data <= 32'h34302578;
         'd5370: data <= 32'h00000a78;         'd5371: data <= 32'h5d64255b;
         'd5372: data <= 32'h6c637263;         'd5373: data <= 32'h20747369;
         'd5374: data <= 32'h20202020;         'd5375: data <= 32'h203a2020;
         'd5376: data <= 32'h30257830;         'd5377: data <= 32'h000a7834;
         'd5378: data <= 32'h5d64255b;         'd5379: data <= 32'h6d637263;
         'd5380: data <= 32'h69727461;         'd5381: data <= 32'h20202078;
         'd5382: data <= 32'h203a2020;         'd5383: data <= 32'h30257830;
         'd5384: data <= 32'h000a7834;         'd5385: data <= 32'h5d64255b;
         'd5386: data <= 32'h73637263;         'd5387: data <= 32'h65746174;
         'd5388: data <= 32'h20202020;         'd5389: data <= 32'h203a2020;
         'd5390: data <= 32'h30257830;         'd5391: data <= 32'h000a7834;
         'd5392: data <= 32'h5d64255b;         'd5393: data <= 32'h66637263;
         'd5394: data <= 32'h6c616e69;         'd5395: data <= 32'h20202020;
         'd5396: data <= 32'h203a2020;         'd5397: data <= 32'h30257830;
         'd5398: data <= 32'h000a7834;         'd5399: data <= 32'h72726f43;
         'd5400: data <= 32'h20746365;         'd5401: data <= 32'h7265706f;
         'd5402: data <= 32'h6f697461;         'd5403: data <= 32'h6176206e;
         'd5404: data <= 32'h6164696c;         'd5405: data <= 32'h2e646574;
         'd5406: data <= 32'h65655320;         'd5407: data <= 32'h41455220;
         'd5408: data <= 32'h2e454d44;         'd5409: data <= 32'h6620646d;
         'd5410: data <= 32'h7220726f;         'd5411: data <= 32'h61206e75;
         'd5412: data <= 32'h7220646e;         'd5413: data <= 32'h726f7065;
         'd5414: data <= 32'h676e6974;         'd5415: data <= 32'h6c757220;
         'd5416: data <= 32'h0a2e7365;         'd5417: data <= 32'h00000000;
         'd5418: data <= 32'h6f727245;         'd5419: data <= 32'h64207372;
         'd5420: data <= 32'h63657465;         'd5421: data <= 32'h0a646574;
         'd5422: data <= 32'h00000000;         'd5423: data <= 32'h6e6e6143;
         'd5424: data <= 32'h7620746f;         'd5425: data <= 32'h64696c61;
         'd5426: data <= 32'h20657461;         'd5427: data <= 32'h7265706f;
         'd5428: data <= 32'h6f697461;         'd5429: data <= 32'h6f66206e;
         'd5430: data <= 32'h68742072;         'd5431: data <= 32'h20657365;
         'd5432: data <= 32'h64656573;         'd5433: data <= 32'h6c617620;
         'd5434: data <= 32'h2c736575;         'd5435: data <= 32'h656c7020;
         'd5436: data <= 32'h20657361;         'd5437: data <= 32'h706d6f63;
         'd5438: data <= 32'h20657261;         'd5439: data <= 32'h68746977;
         'd5440: data <= 32'h73657220;         'd5441: data <= 32'h73746c75;
         'd5442: data <= 32'h206e6f20;         'd5443: data <= 32'h6e6b2061;
         'd5444: data <= 32'h206e776f;         'd5445: data <= 32'h74616c70;
         'd5446: data <= 32'h6d726f66;         'd5447: data <= 32'h00000a2e;
         'd5448: data <= 32'h32313035;         'd5449: data <= 32'h00000000;
         'd5450: data <= 32'h34333231;         'd5451: data <= 32'h00000000;
         'd5452: data <= 32'h3437382d;         'd5453: data <= 32'h00000000;
         'd5454: data <= 32'h3232312b;         'd5455: data <= 32'h00000000;
         'd5456: data <= 32'h352e3533;         'd5457: data <= 32'h30303434;
         'd5458: data <= 32'h00000000;         'd5459: data <= 32'h3332312e;
         'd5460: data <= 32'h30303534;         'd5461: data <= 32'h00000000;
         'd5462: data <= 32'h3031312d;         'd5463: data <= 32'h3030372e;
         'd5464: data <= 32'h00000000;         'd5465: data <= 32'h362e302b;
         'd5466: data <= 32'h30303434;         'd5467: data <= 32'h00000000;
         'd5468: data <= 32'h30352e35;         'd5469: data <= 32'h332b6530;
         'd5470: data <= 32'h00000000;         'd5471: data <= 32'h32312e2d;
         'd5472: data <= 32'h322d6533;         'd5473: data <= 32'h00000000;
         'd5474: data <= 32'h6537382d;         'd5475: data <= 32'h3233382b;
         'd5476: data <= 32'h00000000;         'd5477: data <= 32'h362e302b;
         'd5478: data <= 32'h32312d65;         'd5479: data <= 32'h00000000;
         'd5480: data <= 32'h332e3054;         'd5481: data <= 32'h46312d65;
         'd5482: data <= 32'h00000000;         'd5483: data <= 32'h542e542d;
         'd5484: data <= 32'h71542b2b;         'd5485: data <= 32'h00000000;
         'd5486: data <= 32'h2e335431;         'd5487: data <= 32'h7a346534;
         'd5488: data <= 32'h00000000;         'd5489: data <= 32'h302e3433;
         'd5490: data <= 32'h5e542d65;         'd5491: data <= 32'h00000000;
         'd5492: data <= 32'h800031bc;         'd5493: data <= 32'h80003478;
         'd5494: data <= 32'h8000324c;         'd5495: data <= 32'h80003398;
         'd5496: data <= 32'h800032cc;         'd5497: data <= 32'h8000332c;
         'd5498: data <= 32'h800033f0;         'd5499: data <= 32'h80003444;
         'd5500: data <= 32'h80003550;         'd5501: data <= 32'h80003514;
         'd5502: data <= 32'h80003520;         'd5503: data <= 32'h8000352c;
         'd5504: data <= 32'h80003538;         'd5505: data <= 32'h80003544;
         'd5506: data <= 32'h4f525245;         'd5507: data <= 32'h50203a52;
         'd5508: data <= 32'h7361656c;         'd5509: data <= 32'h6f6d2065;
         'd5510: data <= 32'h79666964;         'd5511: data <= 32'h65687420;
         'd5512: data <= 32'h74616420;         'd5513: data <= 32'h70797461;
         'd5514: data <= 32'h69207365;         'd5515: data <= 32'h6f63206e;
         'd5516: data <= 32'h705f6572;         'd5517: data <= 32'h6d74726f;
         'd5518: data <= 32'h21682e65;         'd5519: data <= 32'h0000000a;
         'd5520: data <= 32'h80004130;         'd5521: data <= 32'h80004178;
         'd5522: data <= 32'h80004178;         'd5523: data <= 32'h80004154;
         'd5524: data <= 32'h80004178;         'd5525: data <= 32'h80004178;
         'd5526: data <= 32'h80004178;         'd5527: data <= 32'h80004178;
         'd5528: data <= 32'h80004178;         'd5529: data <= 32'h80004178;
         'd5530: data <= 32'h80004178;         'd5531: data <= 32'h8000410c;
         'd5532: data <= 32'h80004178;         'd5533: data <= 32'h800040e8;
         'd5534: data <= 32'h80004178;         'd5535: data <= 32'h80004178;
         'd5536: data <= 32'h800040c4;         'd5537: data <= 32'h8000431c;
         'd5538: data <= 32'h800043b4;         'd5539: data <= 32'h8000437c;
         'd5540: data <= 32'h800043b4;         'd5541: data <= 32'h800042d8;
         'd5542: data <= 32'h800043b4;         'd5543: data <= 32'h800043b4;
         'd5544: data <= 32'h800043b4;         'd5545: data <= 32'h800043b4;
         'd5546: data <= 32'h800043b4;         'd5547: data <= 32'h800043b4;
         'd5548: data <= 32'h800043b4;         'd5549: data <= 32'h80004360;
         'd5550: data <= 32'h800043b4;         'd5551: data <= 32'h800043b4;
         'd5552: data <= 32'h800043b4;         'd5553: data <= 32'h800043b4;
         'd5554: data <= 32'h800043b4;         'd5555: data <= 32'h80004398;
         'd5556: data <= 32'h800049dc;         'd5557: data <= 32'h80004a10;
         'd5558: data <= 32'h80004a10;         'd5559: data <= 32'h80004a10;
         'd5560: data <= 32'h80004a10;         'd5561: data <= 32'h80004a10;
         'd5562: data <= 32'h80004a10;         'd5563: data <= 32'h80004a10;
         'd5564: data <= 32'h80004a10;         'd5565: data <= 32'h80004a10;
         'd5566: data <= 32'h80004a10;         'd5567: data <= 32'h80004a10;
         'd5568: data <= 32'h80004a10;         'd5569: data <= 32'h80004a10;
         'd5570: data <= 32'h80004a10;         'd5571: data <= 32'h80004a10;
         'd5572: data <= 32'h80004a10;         'd5573: data <= 32'h80004a10;
         'd5574: data <= 32'h80004a10;         'd5575: data <= 32'h80004a10;
         'd5576: data <= 32'h80004a10;         'd5577: data <= 32'h80004a10;
         'd5578: data <= 32'h80004a10;         'd5579: data <= 32'h80004a10;
         'd5580: data <= 32'h80004a10;         'd5581: data <= 32'h80004a10;
         'd5582: data <= 32'h80004a10;         'd5583: data <= 32'h80004a10;
         'd5584: data <= 32'h80004a10;         'd5585: data <= 32'h80004a10;
         'd5586: data <= 32'h80004a10;         'd5587: data <= 32'h80004a10;
         'd5588: data <= 32'h80004a10;         'd5589: data <= 32'h80004a10;
         'd5590: data <= 32'h80004a10;         'd5591: data <= 32'h80004a10;
         'd5592: data <= 32'h80004a10;         'd5593: data <= 32'h80004a10;
         'd5594: data <= 32'h80004a10;         'd5595: data <= 32'h80004a10;
         'd5596: data <= 32'h80004a10;         'd5597: data <= 32'h80004a10;
         'd5598: data <= 32'h80004a10;         'd5599: data <= 32'h80004a10;
         'd5600: data <= 32'h80004a10;         'd5601: data <= 32'h80004a10;
         'd5602: data <= 32'h80004a10;         'd5603: data <= 32'h80004a10;
         'd5604: data <= 32'h80004a10;         'd5605: data <= 32'h80004a10;
         'd5606: data <= 32'h80004a10;         'd5607: data <= 32'h800043f4;
         'd5608: data <= 32'h80004a10;         'd5609: data <= 32'h80004a10;
         'd5610: data <= 32'h80004a10;         'd5611: data <= 32'h80004a10;
         'd5612: data <= 32'h80004a10;         'd5613: data <= 32'h80004a10;
         'd5614: data <= 32'h80004a10;         'd5615: data <= 32'h80004a10;
         'd5616: data <= 32'h80004a10;         'd5617: data <= 32'h800043f4;
         'd5618: data <= 32'h80004740;         'd5619: data <= 32'h800043f4;
         'd5620: data <= 32'h80004a10;         'd5621: data <= 32'h80004a10;
         'd5622: data <= 32'h80004a10;         'd5623: data <= 32'h80004a10;
         'd5624: data <= 32'h800043f4;         'd5625: data <= 32'h80004a10;
         'd5626: data <= 32'h80004a10;         'd5627: data <= 32'h80004a10;
         'd5628: data <= 32'h80004a10;         'd5629: data <= 32'h80004a10;
         'd5630: data <= 32'h800043f4;         'd5631: data <= 32'h80004970;
         'd5632: data <= 32'h80004a10;         'd5633: data <= 32'h80004a10;
         'd5634: data <= 32'h8000481c;         'd5635: data <= 32'h80004a10;
         'd5636: data <= 32'h800043f4;         'd5637: data <= 32'h80004a10;
         'd5638: data <= 32'h80004a10;         'd5639: data <= 32'h800043f4;
         'd5640: data <= 32'h2d200d0a;         'd5641: data <= 32'h2d2d2d2d;
         'd5642: data <= 32'h2d2d2d2d;         'd5643: data <= 32'h00002d2d;
         'd5644: data <= 32'h43200d0a;         'd5645: data <= 32'h6d65726f;
         'd5646: data <= 32'h206b7261;         'd5647: data <= 32'h72617453;
         'd5648: data <= 32'h00000074;         'd5649: data <= 32'h3340d4b0;
         'd5650: data <= 32'he7146a79;         'd5651: data <= 32'h0000e3c1;
         'd5652: data <= 32'h1199be52;         'd5653: data <= 32'h1fd75608;
         'd5654: data <= 32'h00000747;         'd5655: data <= 32'h39bf5e47;
         'd5656: data <= 32'h8e3ae5a4;         'd5657: data <= 32'h00008d84;
         'd5658: data <= 32'h80005004;         'd5659: data <= 32'h8000500c;
         'd5660: data <= 32'h80005014;         'd5661: data <= 32'h80005520;
         'd5662: data <= 32'h80005528;         'd5663: data <= 32'h80005530;
         'd5664: data <= 32'h80005538;         'd5665: data <= 32'h80005540;
         'd5666: data <= 32'h8000554c;         'd5667: data <= 32'h80005558;
         'd5668: data <= 32'h80005564;         'd5669: data <= 32'h80005570;
         'd5670: data <= 32'h8000557c;         'd5671: data <= 32'h80005588;
         'd5672: data <= 32'h80005594;         'd5673: data <= 32'h800055a0;
         'd5674: data <= 32'h800055ac;         'd5675: data <= 32'h800055b8;
         'd5676: data <= 32'h800055c4;         'd5677: data <= 32'h00000066;
         'd5678: data <= 32'h00000001;
         default: data <= '0;
         endcase
     end
 end
endmodule
